`timescale 1us/1ns





module tbwinequality_red_ts #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000




)();
  reg [FEAT_BITS*FEAT_CNT-1:0] data;
  wire [FEAT_BITS*FEAT_CNT-1:0] testcases [TEST_CNT-1:0];
  reg rst;
  reg clk;
  parameter Nsperiod=50000;
  localparam period=Nsperiod/500;
  localparam halfT=period/2;


assign testcases[0] = 44'h46012229a22;
assign testcases[1] = 44'h58022538633;
assign testcases[2] = 44'h57122338733;
assign testcases[3] = 44'h92912439523;
assign testcases[4] = 44'h46012229a22;
assign testcases[5] = 44'h46012329a22;
assign testcases[6] = 44'h55112337712;
assign testcases[7] = 44'h46001315814;
assign testcases[8] = 44'h55012218823;
assign testcases[9] = 44'h44662459855;
assign testcases[10] = 44'h35112337722;
assign testcases[11] = 44'h44662459855;
assign testcases[12] = 44'h15012335b24;
assign testcases[13] = 44'h555132197c2;
assign testcases[14] = 44'h65334b8a552;
assign testcases[15] = 44'h65334b8a562;
assign testcases[16] = 44'h62912858745;
assign testcases[17] = 44'h5541a338592;
assign testcases[18] = 44'h45142119821;
assign testcases[19] = 44'h52819438472;
assign testcases[20] = 44'h61812638822;
assign testcases[21] = 44'h4352254aa33;
assign testcases[22] = 44'h53313228563;
assign testcases[23] = 44'h64222238522;
assign testcases[24] = 44'h33222528933;
assign testcases[25] = 44'h23312216822;
assign testcases[26] = 44'h43412107723;
assign testcases[27] = 44'h53313228563;
assign testcases[28] = 44'h46012328922;
assign testcases[29] = 44'h56012217823;
assign testcases[30] = 44'h36122447824;
assign testcases[31] = 44'h36022528925;
assign testcases[32] = 44'h56222368533;
assign testcases[33] = 44'h352b294b922;
assign testcases[34] = 44'h12412327822;
assign testcases[35] = 44'h5605211a823;
assign testcases[36] = 44'h55222019936;
assign testcases[37] = 44'h53411318643;
assign testcases[38] = 44'h2b114115a13;
assign testcases[39] = 44'h44652259755;
assign testcases[40] = 44'h44652259755;
assign testcases[41] = 44'h65522429722;
assign testcases[42] = 44'h44329208655;
assign testcases[43] = 44'h56412218785;
assign testcases[44] = 44'h36011107923;
assign testcases[45] = 44'h04211234f2c;
assign testcases[46] = 44'h49713568642;
assign testcases[47] = 44'h62813228623;
assign testcases[48] = 44'h33411107822;
assign testcases[49] = 44'h12612256722;
assign testcases[50] = 44'h66412118542;
assign testcases[51] = 44'h34112216832;
assign testcases[52] = 44'h34111106832;
assign testcases[53] = 44'h63622768622;
assign testcases[54] = 44'h44223746534;
assign testcases[55] = 44'h45132529823;
assign testcases[56] = 44'h83932108433;
assign testcases[57] = 44'h46253b6a742;
assign testcases[58] = 44'h55322439924;
assign testcases[59] = 44'h43522227822;
assign testcases[60] = 44'h63612439932;
assign testcases[61] = 44'h46813468642;
assign testcases[62] = 44'h44312228833;
assign testcases[63] = 44'h37112338823;
assign testcases[64] = 44'h47142107816;
assign testcases[65] = 44'h47142107816;
assign testcases[66] = 44'h44212228923;
assign testcases[67] = 44'h36112117926;
assign testcases[68] = 44'h72912638746;
assign testcases[69] = 44'h56112217865;
assign testcases[70] = 44'h46112318723;
assign testcases[71] = 44'h46412457713;
assign testcases[72] = 44'h46412457713;
assign testcases[73] = 44'h56412229722;
assign testcases[74] = 44'h7292264a753;
assign testcases[75] = 44'h63a1222aa35;
assign testcases[76] = 44'h63a1222aa35;
assign testcases[77] = 44'h37022318a26;
assign testcases[78] = 44'h37212247824;
assign testcases[79] = 44'h56312668582;
assign testcases[80] = 44'h24312017822;
assign testcases[81] = 44'h53b1c539592;
assign testcases[82] = 44'h44812548822;
assign testcases[83] = 44'h4641a338582;
assign testcases[84] = 44'h22812437945;
assign testcases[85] = 44'h35212427824;
assign testcases[86] = 44'h644134782f4;
assign testcases[87] = 44'h44411218833;
assign testcases[88] = 44'h73713779593;
assign testcases[89] = 44'h35112219921;
assign testcases[90] = 44'h54412987623;
assign testcases[91] = 44'h644134782f4;
assign testcases[92] = 44'h645134782f3;
assign testcases[93] = 44'h44411218833;
assign testcases[94] = 44'h1a111944d15;
assign testcases[95] = 44'h05321464e3b;
assign testcases[96] = 44'h37022218926;
assign testcases[97] = 44'h34412017632;
assign testcases[98] = 44'h49122108823;
assign testcases[99] = 44'h55312328721;
assign testcases[100] = 44'h55512228834;
assign testcases[101] = 44'h54512217725;
assign testcases[102] = 44'h55312328721;
assign testcases[103] = 44'h55412238722;
assign testcases[104] = 44'h44412127712;
assign testcases[105] = 44'h55412238722;
assign testcases[106] = 44'h53b1c448492;
assign testcases[107] = 44'h26512338942;
assign testcases[108] = 44'h52822449853;
assign testcases[109] = 44'h57813888632;
assign testcases[110] = 44'h55312227663;
assign testcases[111] = 44'h55112267533;
assign testcases[112] = 44'h55212367533;
assign testcases[113] = 44'h8272252a733;
assign testcases[114] = 44'h55312227663;
assign testcases[115] = 44'h73512338435;
assign testcases[116] = 44'h55412229834;
assign testcases[117] = 44'h55212118822;
assign testcases[118] = 44'h65113337636;
assign testcases[119] = 44'h36112557822;
assign testcases[120] = 44'h4a114257721;
assign testcases[121] = 44'h65113337636;
assign testcases[122] = 44'h46022009922;
assign testcases[123] = 44'h56022229923;
assign testcases[124] = 44'h54312557813;
assign testcases[125] = 44'h6511465a542;
assign testcases[126] = 44'h5d012007a26;
assign testcases[127] = 44'h5d012007a16;
assign testcases[128] = 44'h55311017965;
assign testcases[129] = 44'h23212116922;
assign testcases[130] = 44'h57913778632;
assign testcases[131] = 44'h14121454b3b;
assign testcases[132] = 44'h14121454b3b;
assign testcases[133] = 44'h34011416823;
assign testcases[134] = 44'h5a112317624;
assign testcases[135] = 44'h57212338653;
assign testcases[136] = 44'h57212238643;
assign testcases[137] = 44'h43612328932;
assign testcases[138] = 44'h55312367723;
assign testcases[139] = 44'h55312467723;
assign testcases[140] = 44'h57212338653;
assign testcases[141] = 44'h57212238643;
assign testcases[142] = 44'h12011632c4e;
assign testcases[143] = 44'h23111016822;
assign testcases[144] = 44'h12011632c4e;
assign testcases[145] = 44'h56913788532;
assign testcases[146] = 44'h26012555a24;
assign testcases[147] = 44'h44416258552;
assign testcases[148] = 44'h34222217924;
assign testcases[149] = 44'h53722229a35;
assign testcases[150] = 44'h42812107725;
assign testcases[151] = 44'h74f3f74b0f2;
assign testcases[152] = 44'h45012556824;
assign testcases[153] = 44'h45012556824;
assign testcases[154] = 44'h43752678945;
assign testcases[155] = 44'h43752678945;
assign testcases[156] = 44'h43752678945;
assign testcases[157] = 44'h43752678945;
assign testcases[158] = 44'h46012218922;
assign testcases[159] = 44'h35312458b22;
assign testcases[160] = 44'h49012117623;
assign testcases[161] = 44'h46002218572;
assign testcases[162] = 44'h54112417724;
assign testcases[163] = 44'h4547287a822;
assign testcases[164] = 44'h45472879822;
assign testcases[165] = 44'h56812357633;
assign testcases[166] = 44'h36212456824;
assign testcases[167] = 44'h45012426811;
assign testcases[168] = 44'h36112226925;
assign testcases[169] = 44'h464193373c3;
assign testcases[170] = 44'h58011108802;
assign testcases[171] = 44'h53312118732;
assign testcases[172] = 44'h53312118732;
assign testcases[173] = 44'h45111527928;
assign testcases[174] = 44'h43312127713;
assign testcases[175] = 44'h34112427843;
assign testcases[176] = 44'h43312127713;
assign testcases[177] = 44'h44722228b35;
assign testcases[178] = 44'h38021118923;
assign testcases[179] = 44'h65221228623;
assign testcases[180] = 44'h65221228623;
assign testcases[181] = 44'h65817568572;
assign testcases[182] = 44'h47022328922;
assign testcases[183] = 44'h35312238a22;
assign testcases[184] = 44'h35312238a22;
assign testcases[185] = 44'h62913648723;
assign testcases[186] = 44'h43812338822;
assign testcases[187] = 44'h46222219823;
assign testcases[188] = 44'h54512388623;
assign testcases[189] = 44'h54512488623;
assign testcases[190] = 44'h54622579632;
assign testcases[191] = 44'h33412529a33;
assign testcases[192] = 44'h36232378733;
assign testcases[193] = 44'h45312117723;
assign testcases[194] = 44'h45312117723;
assign testcases[195] = 44'h55512568622;
assign testcases[196] = 44'h45522338924;
assign testcases[197] = 44'ha2a11219564;
assign testcases[198] = 44'h18101353a5b;
assign testcases[199] = 44'h3b111216a17;
assign testcases[200] = 44'h72811218655;
assign testcases[201] = 44'h63812989472;
assign testcases[202] = 44'h34212326843;
assign testcases[203] = 44'h33612327822;
assign testcases[204] = 44'h33612327822;
assign testcases[205] = 44'hc2c2221b646;
assign testcases[206] = 44'hc2c2221b646;
assign testcases[207] = 44'h55512667722;
assign testcases[208] = 44'h54422458632;
assign testcases[209] = 44'h92911119755;
assign testcases[210] = 44'h74a1111775a;
assign testcases[211] = 44'h57422238824;
assign testcases[212] = 44'ha4a11119634;
assign testcases[213] = 44'h55411637714;
assign testcases[214] = 44'h57122229643;
assign testcases[215] = 44'h34851679845;
assign testcases[216] = 44'h66312327526;
assign testcases[217] = 44'h57412228822;
assign testcases[218] = 44'h44312227823;
assign testcases[219] = 44'h54522588733;
assign testcases[220] = 44'h52612537822;
assign testcases[221] = 44'h44412347522;
assign testcases[222] = 44'h35111106933;
assign testcases[223] = 44'h66412219734;
assign testcases[224] = 44'h56612339725;
assign testcases[225] = 44'h43422637825;
assign testcases[226] = 44'h658196474c3;
assign testcases[227] = 44'h6822221a833;
assign testcases[228] = 44'h43422637825;
assign testcases[229] = 44'h34422228926;
assign testcases[230] = 44'h14111463a39;
assign testcases[231] = 44'h53112227824;
assign testcases[232] = 44'h63322439843;
assign testcases[233] = 44'h34422228926;
assign testcases[234] = 44'h5a121128721;
assign testcases[235] = 44'h46012328821;
assign testcases[236] = 44'h46012328821;
assign testcases[237] = 44'h46012328822;
assign testcases[238] = 44'h46012328821;
assign testcases[239] = 44'h5a121128721;
assign testcases[240] = 44'h66617138372;
assign testcases[241] = 44'ha391211b546;
assign testcases[242] = 44'h45212667423;
assign testcases[243] = 44'hf171221c452;
assign testcases[244] = 44'hf171221c452;
assign testcases[245] = 44'h4601211ab64;
assign testcases[246] = 44'h46112338823;
assign testcases[247] = 44'h55322247612;
assign testcases[248] = 44'h44112227813;
assign testcases[249] = 44'h4601211ab64;
assign testcases[250] = 44'h9271132a644;
assign testcases[251] = 44'h45012328944;
assign testcases[252] = 44'h9382211a525;
assign testcases[253] = 44'h47712257623;
assign testcases[254] = 44'h45012328944;
assign testcases[255] = 44'h55432468722;
assign testcases[256] = 44'h72612109632;
assign testcases[257] = 44'h36012238932;
assign testcases[258] = 44'h43c1f228492;
assign testcases[259] = 44'h8282232b855;
assign testcases[260] = 44'h52412427732;
assign testcases[261] = 44'h39112237832;
assign testcases[262] = 44'h54012227824;
assign testcases[263] = 44'h53412527732;
assign testcases[264] = 44'hb582111c456;
assign testcases[265] = 44'ha2812108644;
assign testcases[266] = 44'h5803263cb43;
assign testcases[267] = 44'h5373232885b;
assign testcases[268] = 44'h3512211ac62;
assign testcases[269] = 44'ha183211b764;
assign testcases[270] = 44'h55132638836;
assign testcases[271] = 44'ha183211b764;
assign testcases[272] = 44'h9393243b644;
assign testcases[273] = 44'h57322229732;
assign testcases[274] = 44'h4637265b842;
assign testcases[275] = 44'h55132638836;
assign testcases[276] = 44'h3512211ac62;
assign testcases[277] = 44'ha183211b764;
assign testcases[278] = 44'h8276210965a;
assign testcases[279] = 44'h6355222b845;
assign testcases[280] = 44'ha273211a552;
assign testcases[281] = 44'h42b39108674;
assign testcases[282] = 44'h44221238822;
assign testcases[283] = 44'h6355222b845;
assign testcases[284] = 44'h8513274c743;
assign testcases[285] = 44'h8513274c743;
assign testcases[286] = 44'ha491252b545;
assign testcases[287] = 44'h43222638845;
assign testcases[288] = 44'h64122429855;
assign testcases[289] = 44'ha383275d662;
assign testcases[290] = 44'h64122429855;
assign testcases[291] = 44'h91819119745;
assign testcases[292] = 44'h8542242b635;
assign testcases[293] = 44'h33422117834;
assign testcases[294] = 44'hc283243d453;
assign testcases[295] = 44'h9472211c433;
assign testcases[296] = 44'h88622649524;
assign testcases[297] = 44'h4611221ac43;
assign testcases[298] = 44'h4602211bc53;
assign testcases[299] = 44'h3611222ac43;
assign testcases[300] = 44'h44122428826;
assign testcases[301] = 44'h91811118634;
assign testcases[302] = 44'h5622221ba44;
assign testcases[303] = 44'h46215117823;
assign testcases[304] = 44'h56a13258622;
assign testcases[305] = 44'h8482111b522;
assign testcases[306] = 44'h45512138822;
assign testcases[307] = 44'h8372510b633;
assign testcases[308] = 44'h8372510b633;
assign testcases[309] = 44'h42611218823;
assign testcases[310] = 44'h8482111b522;
assign testcases[311] = 44'h54412367722;
assign testcases[312] = 44'h64522459733;
assign testcases[313] = 44'h64522779722;
assign testcases[314] = 44'h43522647836;
assign testcases[315] = 44'h43522437936;
assign testcases[316] = 44'h7543285b734;
assign testcases[317] = 44'h7722274a735;
assign testcases[318] = 44'h7663253a848;
assign testcases[319] = 44'h7722274a735;
assign testcases[320] = 44'h7663253a848;
assign testcases[321] = 44'h7543255b633;
assign testcases[322] = 44'h55122119732;
assign testcases[323] = 44'h8572284a743;
assign testcases[324] = 44'h843b232d532;
assign testcases[325] = 44'h843b232d532;
assign testcases[326] = 44'ha4b33109448;
assign testcases[327] = 44'h84843109758;
assign testcases[328] = 44'hc2a2211c533;
assign testcases[329] = 44'h94611119633;
assign testcases[330] = 44'h83a2322963a;
assign testcases[331] = 44'h83a2322963a;
assign testcases[332] = 44'h55431568622;
assign testcases[333] = 44'h55112327526;
assign testcases[334] = 44'h56022427848;
assign testcases[335] = 44'ha683311b559;
assign testcases[336] = 44'h6371111684a;
assign testcases[337] = 44'h53522639735;
assign testcases[338] = 44'hb492265d568;
assign testcases[339] = 44'hb292221b5a3;
assign testcases[340] = 44'hb282121c582;
assign testcases[341] = 44'h83821118657;
assign testcases[342] = 44'h9381310a743;
assign testcases[343] = 44'h9381310a743;
assign testcases[344] = 44'ha582211c546;
assign testcases[345] = 44'h36011939b54;
assign testcases[346] = 44'h38022426b5a;
assign testcases[347] = 44'hd4b2211a469;
assign testcases[348] = 44'h75522329564;
assign testcases[349] = 44'h6702221b852;
assign testcases[350] = 44'h9642342c764;
assign testcases[351] = 44'h6702221b852;
assign testcases[352] = 44'h46022219742;
assign testcases[353] = 44'hd4d4354e64b;
assign testcases[354] = 44'h21611991629;
assign testcases[355] = 44'h37022416a3b;
assign testcases[356] = 44'ha382263c756;
assign testcases[357] = 44'h83b23218648;
assign testcases[358] = 44'ha3b2321c555;
assign testcases[359] = 44'hb3b2222d533;
assign testcases[360] = 44'h56412348642;
assign testcases[361] = 44'h6452252a864;
assign testcases[362] = 44'ha5b2212b424;
assign testcases[363] = 44'hb4a1211a354;
assign testcases[364] = 44'hc5b5212e444;
assign testcases[365] = 44'h83833119768;
assign testcases[366] = 44'hc5b5212e444;
assign testcases[367] = 44'h85a2221c531;
assign testcases[368] = 44'h8282434b632;
assign testcases[369] = 44'h72822117689;
assign testcases[370] = 44'h37021839a44;
assign testcases[371] = 44'h51611218751;
assign testcases[372] = 44'h62811628775;
assign testcases[373] = 44'h45413247432;
assign testcases[374] = 44'hd3a3212d356;
assign testcases[375] = 44'ha5b4311a358;
assign testcases[376] = 44'ha482242c776;
assign testcases[377] = 44'h72822117689;
assign testcases[378] = 44'ha6b6211a56c;
assign testcases[379] = 44'h53622539746;
assign testcases[380] = 44'h52712219652;
assign testcases[381] = 44'hd3b2242d454;
assign testcases[382] = 44'h52712219652;
assign testcases[383] = 44'h52712219652;
assign testcases[384] = 44'h44412539942;
assign testcases[385] = 44'h46122229943;
assign testcases[386] = 44'h55412529842;
assign testcases[387] = 44'h56212428723;
assign testcases[388] = 44'h54412539942;
assign testcases[389] = 44'h7352232a644;
assign testcases[390] = 44'h18111253a5b;
assign testcases[391] = 44'hd3b2242d454;
assign testcases[392] = 44'h73812119623;
assign testcases[393] = 44'h56a13358522;
assign testcases[394] = 44'hb5a2111b424;
assign testcases[395] = 44'ha3c4112c63b;
assign testcases[396] = 44'h37083f7b924;
assign testcases[397] = 44'ha592232a636;
assign testcases[398] = 44'ha592232a636;
assign testcases[399] = 44'h67421227522;
assign testcases[400] = 44'h37083f7b924;
assign testcases[401] = 44'h42511426716;
assign testcases[402] = 44'hb492243c535;
assign testcases[403] = 44'ha582222b535;
assign testcases[404] = 44'h46122319732;
assign testcases[405] = 44'h62711218844;
assign testcases[406] = 44'h74821219636;
assign testcases[407] = 44'ha3b2221b636;
assign testcases[408] = 44'h82934118647;
assign testcases[409] = 44'hb4842629423;
assign testcases[410] = 44'h6352265a833;
assign testcases[411] = 44'h6462254a833;
assign testcases[412] = 44'h47312348732;
assign testcases[413] = 44'h8386211a758;
assign testcases[414] = 44'h6452257a733;
assign testcases[415] = 44'h6746377d772;
assign testcases[416] = 44'h84a13118738;
assign testcases[417] = 44'h35212776915;
assign testcases[418] = 44'ha381311b645;
assign testcases[419] = 44'h37011739b34;
assign testcases[420] = 44'h75522838748;
assign testcases[421] = 44'h38021726a2a;
assign testcases[422] = 44'h49311336816;
assign testcases[423] = 44'h81811119556;
assign testcases[424] = 44'h49311336816;
assign testcases[425] = 44'h38021726a2a;
assign testcases[426] = 44'h36111426927;
assign testcases[427] = 44'h7741211a725;
assign testcases[428] = 44'h64502219632;
assign testcases[429] = 44'hc8a2232b535;
assign testcases[430] = 44'h81811119556;
assign testcases[431] = 44'h55612539622;
assign testcases[432] = 44'ha3b2221733b;
assign testcases[433] = 44'hb3a2211c523;
assign testcases[434] = 44'h8393253b554;
assign testcases[435] = 44'hb3a2211c523;
assign testcases[436] = 44'h56511837724;
assign testcases[437] = 44'h94c3111a537;
assign testcases[438] = 44'h8393253b554;
assign testcases[439] = 44'h35311126432;
assign testcases[440] = 44'hb2c1211a253;
assign testcases[441] = 44'ha3a1111a437;
assign testcases[442] = 44'hf6c3212f337;
assign testcases[443] = 44'h84822217638;
assign testcases[444] = 44'h15011114a5a;
assign testcases[445] = 44'h7721211a624;
assign testcases[446] = 44'hb3a2274b545;
assign testcases[447] = 44'h74513118647;
assign testcases[448] = 44'h64412118624;
assign testcases[449] = 44'ha3b2242b536;
assign testcases[450] = 44'ha3b2242b536;
assign testcases[451] = 44'h5381b219472;
assign testcases[452] = 44'h35012428934;
assign testcases[453] = 44'h82a2211b747;
assign testcases[454] = 44'h31611536a37;
assign testcases[455] = 44'h95b5211a63c;
assign testcases[456] = 44'h6562211a825;
assign testcases[457] = 44'h7632263a723;
assign testcases[458] = 44'h82a2211b747;
assign testcases[459] = 44'ha5b1222d621;
assign testcases[460] = 44'h73822319837;
assign testcases[461] = 44'h5542211a732;
assign testcases[462] = 44'h92b22218638;
assign testcases[463] = 44'h56b12578421;
assign testcases[464] = 44'ha291211a342;
assign testcases[465] = 44'h8262221c963;
assign testcases[466] = 44'h8471253a548;
assign testcases[467] = 44'h6472111574e;
assign testcases[468] = 44'ha3b1211c532;
assign testcases[469] = 44'h68002826623;
assign testcases[470] = 44'hc2a2232b435;
assign testcases[471] = 44'h75722538647;
assign testcases[472] = 44'hb392254b555;
assign testcases[473] = 44'h83911108745;
assign testcases[474] = 44'h8281221a652;
assign testcases[475] = 44'h7641211a534;
assign testcases[476] = 44'h72712119743;
assign testcases[477] = 44'h81812119676;
assign testcases[478] = 44'h7641211a534;
assign testcases[479] = 44'h7622211a644;
assign testcases[480] = 44'h826f211f532;
assign testcases[481] = 44'h72922117568;
assign testcases[482] = 44'h8391411a472;
assign testcases[483] = 44'h83a1411a472;
assign testcases[484] = 44'h84b4311843c;
assign testcases[485] = 44'h86611119514;
assign testcases[486] = 44'h86611119514;
assign testcases[487] = 44'h8661110a514;
assign testcases[488] = 44'ha292283c766;
assign testcases[489] = 44'h7362221a844;
assign testcases[490] = 44'h7742253a735;
assign testcases[491] = 44'h7382121684c;
assign testcases[492] = 44'h6382131675c;
assign testcases[493] = 44'h6652254c948;
assign testcases[494] = 44'h33481656929;
assign testcases[495] = 44'h93822118536;
assign testcases[496] = 44'h5441232a931;
assign testcases[497] = 44'h42522968747;
assign testcases[498] = 44'h93822118536;
assign testcases[499] = 44'h6652254c948;
assign testcases[500] = 44'h5441232a931;
assign testcases[501] = 44'h84c6284a559;
assign testcases[502] = 44'h84c6284a559;
assign testcases[503] = 44'h82812119676;
assign testcases[504] = 44'h81712119676;
assign testcases[505] = 44'h84a2221854a;
assign testcases[506] = 44'h81712119676;
assign testcases[507] = 44'h9692210c543;
assign testcases[508] = 44'h8551263b634;
assign testcases[509] = 44'hc2c2252a437;
assign testcases[510] = 44'hb3842429433;
assign testcases[511] = 44'h8551263b634;
assign testcases[512] = 44'h93813329453;
assign testcases[513] = 44'h84a23118438;
assign testcases[514] = 44'h84a23118438;
assign testcases[515] = 44'h6686378d782;
assign testcases[516] = 44'hb584210d649;
assign testcases[517] = 44'h8581511b530;
assign testcases[518] = 44'h91822218638;
assign testcases[519] = 44'h43822968846;
assign testcases[520] = 44'h7182232a954;
assign testcases[521] = 44'h43812329932;
assign testcases[522] = 44'h53822a79863;
assign testcases[523] = 44'h73822889622;
assign testcases[524] = 44'h73822569633;
assign testcases[525] = 44'h8642263b634;
assign testcases[526] = 44'h43822968846;
assign testcases[527] = 44'h33822747847;
assign testcases[528] = 44'h5382273a841;
assign testcases[529] = 44'h86422129422;
assign testcases[530] = 44'h6141201a855;
assign testcases[531] = 44'ha382222c535;
assign testcases[532] = 44'ha382222c535;
assign testcases[533] = 44'h8241232663b;
assign testcases[534] = 44'h8442231c724;
assign testcases[535] = 44'h6141201a855;
assign testcases[536] = 44'h86422129422;
assign testcases[537] = 44'h58412108846;
assign testcases[538] = 44'hc385112d639;
assign testcases[539] = 44'h94c5211b637;
assign testcases[540] = 44'h7543242a733;
assign testcases[541] = 44'h7486111a646;
assign testcases[542] = 44'h77412118524;
assign testcases[543] = 44'h9642233b446;
assign testcases[544] = 44'he2c1211d240;
assign testcases[545] = 44'h6482286a422;
assign testcases[546] = 44'h4541221a943;
assign testcases[547] = 44'h8282111a756;
assign testcases[548] = 44'hb382264b545;
assign testcases[549] = 44'h64814119732;
assign testcases[550] = 44'h34012217723;
assign testcases[551] = 44'h73422329644;
assign testcases[552] = 44'h74422329544;
assign testcases[553] = 44'h1a411754d38;
assign testcases[554] = 44'hf684221f247;
assign testcases[555] = 44'hf684221f247;
assign testcases[556] = 44'h9484321c428;
assign testcases[557] = 44'hf684221f247;
assign testcases[558] = 44'h9484321c428;
assign testcases[559] = 44'hc484212e73b;
assign testcases[560] = 44'hb582211b527;
assign testcases[561] = 44'h64822679622;
assign testcases[562] = 44'h6582296a432;
assign testcases[563] = 44'h42822538734;
assign testcases[564] = 44'hc484212e73b;
assign testcases[565] = 44'hb582211b527;
assign testcases[566] = 44'h6642611b731;
assign testcases[567] = 44'h6642611b731;
assign testcases[568] = 44'h7482611a746;
assign testcases[569] = 44'h23412425a28;
assign testcases[570] = 44'ha383222c766;
assign testcases[571] = 44'h23412425a28;
assign testcases[572] = 44'h81822219535;
assign testcases[573] = 44'h8581232b723;
assign testcases[574] = 44'h8283244b644;
assign testcases[575] = 44'hb282262b654;
assign testcases[576] = 44'h84422109824;
assign testcases[577] = 44'h6482246a733;
assign testcases[578] = 44'h6482246a733;
assign testcases[579] = 44'h82811429523;
assign testcases[580] = 44'hb481210c613;
assign testcases[581] = 44'hb481210c613;
assign testcases[582] = 44'ha481211c612;
assign testcases[583] = 44'ha2812219334;
assign testcases[584] = 44'ha2832c4c746;
assign testcases[585] = 44'h44422229933;
assign testcases[586] = 44'h9282232a575;
assign testcases[587] = 44'h47413458722;
assign testcases[588] = 44'h13411422c4e;
assign testcases[589] = 44'h82821109445;
assign testcases[590] = 44'h6482254a823;
assign testcases[591] = 44'h33812583528;
assign testcases[592] = 44'h6482254a823;
assign testcases[593] = 44'h8493222c721;
assign testcases[594] = 44'h57322429823;
assign testcases[595] = 44'h6578276b722;
assign testcases[596] = 44'hb381111b432;
assign testcases[597] = 44'ha5912119434;
assign testcases[598] = 44'h65312118613;
assign testcases[599] = 44'hb572221c342;
assign testcases[600] = 44'h59412117714;
assign testcases[601] = 44'hc481222c521;
assign testcases[602] = 44'h48022109722;
assign testcases[603] = 44'hc481222c521;
assign testcases[604] = 44'h5522233a532;
assign testcases[605] = 44'h5522211a722;
assign testcases[606] = 44'h73842218849;
assign testcases[607] = 44'h6473263a725;
assign testcases[608] = 44'h8665323f735;
assign testcases[609] = 44'h23332326a2b;
assign testcases[610] = 44'h6192253a822;
assign testcases[611] = 44'hc392211c322;
assign testcases[612] = 44'h46022418734;
assign testcases[613] = 44'h53611217743;
assign testcases[614] = 44'h773142582a4;
assign testcases[615] = 44'h7582264ba23;
assign testcases[616] = 44'h7582264ba23;
assign testcases[617] = 44'ha281231a463;
assign testcases[618] = 44'ha482311c544;
assign testcases[619] = 44'h9372211a452;
assign testcases[620] = 44'h55432369732;
assign testcases[621] = 44'h55432369732;
assign testcases[622] = 44'h85412219523;
assign testcases[623] = 44'h54422529969;
assign testcases[624] = 44'h3605353b944;
assign testcases[625] = 44'h3605353b944;
assign testcases[626] = 44'h6551211a822;
assign testcases[627] = 44'h6551211a822;
assign testcases[628] = 44'h65422119732;
assign testcases[629] = 44'h46423447632;
assign testcases[630] = 44'h65422119732;
assign testcases[631] = 44'h8292211a633;
assign testcases[632] = 44'h43222527725;
assign testcases[633] = 44'h8943225d937;
assign testcases[634] = 44'h53312a57723;
assign testcases[635] = 44'h68011526723;
assign testcases[636] = 44'h78422789622;
assign testcases[637] = 44'h78422789622;
assign testcases[638] = 44'h49213117834;
assign testcases[639] = 44'h626115386a5;
assign testcases[640] = 44'h8572232b832;
assign testcases[641] = 44'h7572254b933;
assign testcases[642] = 44'h8572232b832;
assign testcases[643] = 44'h7572254b933;
assign testcases[644] = 44'h8572232b832;
assign testcases[645] = 44'h5626310a834;
assign testcases[646] = 44'h46133118834;
assign testcases[647] = 44'h58012108726;
assign testcases[648] = 44'h64521217737;
assign testcases[649] = 44'h33481586527;
assign testcases[650] = 44'h9361321a223;
assign testcases[651] = 44'h7842288d837;
assign testcases[652] = 44'hf3a7254935f;
assign testcases[653] = 44'h72922219529;
assign testcases[654] = 44'h64822119413;
assign testcases[655] = 44'h7532243c532;
assign testcases[656] = 44'h9361321a223;
assign testcases[657] = 44'ha4912529235;
assign testcases[658] = 44'h44112118753;
assign testcases[659] = 44'h48042108826;
assign testcases[660] = 44'h44112118753;
assign testcases[661] = 44'h43512329731;
assign testcases[662] = 44'h45112218843;
assign testcases[663] = 44'h82711109444;
assign testcases[664] = 44'hb381233c434;
assign testcases[665] = 44'h75212529523;
assign testcases[666] = 44'h54616119633;
assign testcases[667] = 44'h9271211a332;
assign testcases[668] = 44'h87721318526;
assign testcases[669] = 44'h9271211a332;
assign testcases[670] = 44'h33422727724;
assign testcases[671] = 44'h57312108623;
assign testcases[672] = 44'h7c512789523;
assign testcases[673] = 44'h57312108623;
assign testcases[674] = 44'h9371211a432;
assign testcases[675] = 44'h7361121a734;
assign testcases[676] = 44'h9371211a432;
assign testcases[677] = 44'h67222219814;
assign testcases[678] = 44'h57222a5a924;
assign testcases[679] = 44'h92731428523;
assign testcases[680] = 44'hc391232c421;
assign testcases[681] = 44'h54412317624;
assign testcases[682] = 44'h64512739723;
assign testcases[683] = 44'h57421118827;
assign testcases[684] = 44'h79522889612;
assign testcases[685] = 44'h57421118827;
assign testcases[686] = 44'h46312328932;
assign testcases[687] = 44'h6642232b723;
assign testcases[688] = 44'h46111107812;
assign testcases[689] = 44'h53814119772;
assign testcases[690] = 44'h4c042108b26;
assign testcases[691] = 44'h7942225b923;
assign testcases[692] = 44'h6481b339481;
assign testcases[693] = 44'h6452257a732;
assign testcases[694] = 44'h6452257a732;
assign testcases[695] = 44'h14001422f3b;
assign testcases[696] = 44'h36011218933;
assign testcases[697] = 44'h36011218933;
assign testcases[698] = 44'h7543244c723;
assign testcases[699] = 44'ha391211a536;
assign testcases[700] = 44'h8a72265a424;
assign testcases[701] = 44'h36011218933;
assign testcases[702] = 44'h36011218932;
assign testcases[703] = 44'h43822548743;
assign testcases[704] = 44'h67112109723;
assign testcases[705] = 44'h5a26223a824;
assign testcases[706] = 44'h37112216814;
assign testcases[707] = 44'h44322328825;
assign testcases[708] = 44'h55221227838;
assign testcases[709] = 44'h7281132a734;
assign testcases[710] = 44'h8a72254a424;
assign testcases[711] = 44'h6552236b833;
assign testcases[712] = 44'h6603232b812;
assign testcases[713] = 44'h53622229812;
assign testcases[714] = 44'h87422549723;
assign testcases[715] = 44'h44322328712;
assign testcases[716] = 44'h53622229812;
assign testcases[717] = 44'h44222228624;
assign testcases[718] = 44'h55112219613;
assign testcases[719] = 44'h46032429923;
assign testcases[720] = 44'h55112219613;
assign testcases[721] = 44'h6442286a522;
assign testcases[722] = 44'h43122328624;
assign testcases[723] = 44'h425118783c3;
assign testcases[724] = 44'h4b222107a37;
assign testcases[725] = 44'h66322109725;
assign testcases[726] = 44'h5712242b947;
assign testcases[727] = 44'h35011108933;
assign testcases[728] = 44'h35011108933;
assign testcases[729] = 44'h38032636b2b;
assign testcases[730] = 44'h75b2a22a533;
assign testcases[731] = 44'h6823210b928;
assign testcases[732] = 44'h48012218813;
assign testcases[733] = 44'h34522349a33;
assign testcases[734] = 44'h4531222a932;
assign testcases[735] = 44'h49213217723;
assign testcases[736] = 44'h49213217723;
assign testcases[737] = 44'h5502243ca32;
assign testcases[738] = 44'h6442266a522;
assign testcases[739] = 44'h6602242a832;
assign testcases[740] = 44'h57542218938;
assign testcases[741] = 44'h74422689623;
assign testcases[742] = 44'h35011218932;
assign testcases[743] = 44'ha392255c524;
assign testcases[744] = 44'h9392255c523;
assign testcases[745] = 44'h44312219a43;
assign testcases[746] = 44'h52622239711;
assign testcases[747] = 44'h62622349712;
assign testcases[748] = 44'h44312219a43;
assign testcases[749] = 44'h44312219a43;
assign testcases[750] = 44'h56222429723;
assign testcases[751] = 44'h56222429723;
assign testcases[752] = 44'h45222539832;
assign testcases[753] = 44'h56222429723;
assign testcases[754] = 44'h54b1b318472;
assign testcases[755] = 44'h59111526a16;
assign testcases[756] = 44'h29011326b17;
assign testcases[757] = 44'h58012218623;
assign testcases[758] = 44'h58012218623;
assign testcases[759] = 44'h6332275a622;
assign testcases[760] = 44'h65422269623;
assign testcases[761] = 44'h76412129613;
assign testcases[762] = 44'h66012218724;
assign testcases[763] = 44'h76412129613;
assign testcases[764] = 44'h6622222a723;
assign testcases[765] = 44'h7622222a723;
assign testcases[766] = 44'h65322249522;
assign testcases[767] = 44'h4552235b933;
assign testcases[768] = 44'h45022559a23;
assign testcases[769] = 44'h57012118823;
assign testcases[770] = 44'h45022559a23;
assign testcases[771] = 44'h76422589722;
assign testcases[772] = 44'h75422589722;
assign testcases[773] = 44'h53514028763;
assign testcases[774] = 44'h53514028763;
assign testcases[775] = 44'h4a022117914;
assign testcases[776] = 44'h37326127835;
assign testcases[777] = 44'h36326117825;
assign testcases[778] = 44'h53532129835;
assign testcases[779] = 44'h44022559a33;
assign testcases[780] = 44'h35015228732;
assign testcases[781] = 44'h34223229c33;
assign testcases[782] = 44'h68122659824;
assign testcases[783] = 44'h34223229c33;
assign testcases[784] = 44'h45022449a23;
assign testcases[785] = 44'h8372223a623;
assign testcases[786] = 44'h8372223a623;
assign testcases[787] = 44'h8541243b624;
assign testcases[788] = 44'h8541243b624;
assign testcases[789] = 44'h66322569422;
assign testcases[790] = 44'h43722448733;
assign testcases[791] = 44'h6632257a623;
assign testcases[792] = 44'h45022459933;
assign testcases[793] = 44'h45021107826;
assign testcases[794] = 44'h8292111652a;
assign testcases[795] = 44'h98523139384;
assign testcases[796] = 44'h64523539543;
assign testcases[797] = 44'h73711526656;
assign testcases[798] = 44'h7453210a726;
assign testcases[799] = 44'h7453210a726;
assign testcases[800] = 44'h45132667622;
assign testcases[801] = 44'h65131219614;
assign testcases[802] = 44'h15011353a6b;
assign testcases[803] = 44'h45123328633;
assign testcases[804] = 44'h54422118724;
assign testcases[805] = 44'h5262110474b;
assign testcases[806] = 44'h5161110474a;
assign testcases[807] = 44'h5262110474b;
assign testcases[808] = 44'h44214108752;
assign testcases[809] = 44'h44522118625;
assign testcases[810] = 44'h44221107715;
assign testcases[811] = 44'hc492211c436;
assign testcases[812] = 44'h9452242a646;
assign testcases[813] = 44'h33412105927;
assign testcases[814] = 44'hb392242b647;
assign testcases[815] = 44'h9452242a646;
assign testcases[816] = 44'h7433221a625;
assign testcases[817] = 44'h92712416749;
assign testcases[818] = 44'h47022527712;
assign testcases[819] = 44'h6623223b723;
assign testcases[820] = 44'h36012217833;
assign testcases[821] = 44'h03011322c4e;
assign testcases[822] = 44'h35212328b33;
assign testcases[823] = 44'h35212328b33;
assign testcases[824] = 44'h44421118625;
assign testcases[825] = 44'h44222327826;
assign testcases[826] = 44'h42521106836;
assign testcases[827] = 44'h44222327826;
assign testcases[828] = 44'h5512172594b;
assign testcases[829] = 44'h25112314a47;
assign testcases[830] = 44'h46121107826;
assign testcases[831] = 44'h25112314a47;
assign testcases[832] = 44'h8471472a854;
assign testcases[833] = 44'ha471483a854;
assign testcases[834] = 44'h66412318712;
assign testcases[835] = 44'h46211638822;
assign testcases[836] = 44'h32420851718;
assign testcases[837] = 44'h32420851718;
assign testcases[838] = 44'h82612218657;
assign testcases[839] = 44'h24112318914;
assign testcases[840] = 44'h93822229649;
assign testcases[841] = 44'h36023517935;
assign testcases[842] = 44'h84723748646;
assign testcases[843] = 44'h46612257732;
assign testcases[844] = 44'h81711627655;
assign testcases[845] = 44'h36312318b33;
assign testcases[846] = 44'h36312318b33;
assign testcases[847] = 44'h46312229a44;
assign testcases[848] = 44'h36312318b33;
assign testcases[849] = 44'h36312218b33;
assign testcases[850] = 44'h73712218723;
assign testcases[851] = 44'h73712218723;
assign testcases[852] = 44'h53522679673;
assign testcases[853] = 44'h73612938946;
assign testcases[854] = 44'h73612938946;
assign testcases[855] = 44'h47022206a48;
assign testcases[856] = 44'h73612938946;
assign testcases[857] = 44'h52522327847;
assign testcases[858] = 44'ha2811418535;
assign testcases[859] = 44'h35412315857;
assign testcases[860] = 44'h45122349a23;
assign testcases[861] = 44'h2ab11354c38;
assign testcases[862] = 44'h43521117615;
assign testcases[863] = 44'h45122449a23;
assign testcases[864] = 44'h45122349a23;
assign testcases[865] = 44'h46122359a23;
assign testcases[866] = 44'h34422315857;
assign testcases[867] = 44'h34412315857;
assign testcases[868] = 44'h35412315857;
assign testcases[869] = 44'h46012627936;
assign testcases[870] = 44'h47011724828;
assign testcases[871] = 44'h35012826a25;
assign testcases[872] = 44'h43411627924;
assign testcases[873] = 44'h61611106627;
assign testcases[874] = 44'h83712108538;
assign testcases[875] = 44'h62623117748;
assign testcases[876] = 44'h44011106826;
assign testcases[877] = 44'h47011724828;
assign testcases[878] = 44'h65332749624;
assign testcases[879] = 44'h45122459a23;
assign testcases[880] = 44'h75312217524;
assign testcases[881] = 44'h47011726937;
assign testcases[882] = 44'h52525316649;
assign testcases[883] = 44'h45122459a23;
assign testcases[884] = 44'h65332749624;
assign testcases[885] = 44'h6722221a835;
assign testcases[886] = 44'h6722221a735;
assign testcases[887] = 44'h94621637549;
assign testcases[888] = 44'h35022736927;
assign testcases[889] = 44'h9956355f632;
assign testcases[890] = 44'h42412737924;
assign testcases[891] = 44'h46022359a23;
assign testcases[892] = 44'h84412219632;
assign testcases[893] = 44'h46022359a23;
assign testcases[894] = 44'h46012459a23;
assign testcases[895] = 44'h45022626926;
assign testcases[896] = 44'h5262242574a;
assign testcases[897] = 44'h45022626926;
assign testcases[898] = 44'h5262242574a;
assign testcases[899] = 44'h5a03210a926;
assign testcases[900] = 44'h62621227838;
assign testcases[901] = 44'h46222329b36;
assign testcases[902] = 44'h46222329b36;
assign testcases[903] = 44'h35161217826;
assign testcases[904] = 44'h35161217826;
assign testcases[905] = 44'h75322369623;
assign testcases[906] = 44'h45422247846;
assign testcases[907] = 44'h25012106b28;
assign testcases[908] = 44'h44222736926;
assign testcases[909] = 44'h42601104728;
assign testcases[910] = 44'h7383300762c;
assign testcases[911] = 44'h6279300b636;
assign testcases[912] = 44'h84721108739;
assign testcases[913] = 44'h73742007739;
assign testcases[914] = 44'h42601104728;
assign testcases[915] = 44'h62612006739;
assign testcases[916] = 44'h17314135b36;
assign testcases[917] = 44'h3359262a834;
assign testcases[918] = 44'h53512747746;
assign testcases[919] = 44'h55212826858;
assign testcases[920] = 44'h73622219625;
assign testcases[921] = 44'h53512747746;
assign testcases[922] = 44'h55212826858;
assign testcases[923] = 44'h3359262a834;
assign testcases[924] = 44'h64421316657;
assign testcases[925] = 44'h61611c47956;
assign testcases[926] = 44'h71521b49954;
assign testcases[927] = 44'h56312249622;
assign testcases[928] = 44'h64421316657;
assign testcases[929] = 44'h62631215749;
assign testcases[930] = 44'h35012219c45;
assign testcases[931] = 44'h45012329933;
assign testcases[932] = 44'h43512638923;
assign testcases[933] = 44'h45012329933;
assign testcases[934] = 44'h35012219c45;
assign testcases[935] = 44'h62621446848;
assign testcases[936] = 44'h62621446848;
assign testcases[937] = 44'ha6812119435;
assign testcases[938] = 44'h4362152484b;
assign testcases[939] = 44'h24312105b27;
assign testcases[940] = 44'h7281231684a;
assign testcases[941] = 44'h8284221662a;
assign testcases[942] = 44'h8362233a634;
assign testcases[943] = 44'h7452222a633;
assign testcases[944] = 44'h52832216739;
assign testcases[945] = 44'h84712117547;
assign testcases[946] = 44'h84942219769;
assign testcases[947] = 44'h5281210573a;
assign testcases[948] = 44'h60712216849;
assign testcases[949] = 44'h60712216849;
assign testcases[950] = 44'h60712216849;
assign testcases[951] = 44'h5281210573a;
assign testcases[952] = 44'h52611106737;
assign testcases[953] = 44'h82811105639;
assign testcases[954] = 44'h43622106929;
assign testcases[955] = 44'h61812218835;
assign testcases[956] = 44'h63813107737;
assign testcases[957] = 44'h73812237727;
assign testcases[958] = 44'h35223526947;
assign testcases[959] = 44'h55112219834;
assign testcases[960] = 44'h64411426557;
assign testcases[961] = 44'h45212117732;
assign testcases[962] = 44'h35013118833;
assign testcases[963] = 44'h62612416537;
assign testcases[964] = 44'h64411426557;
assign testcases[965] = 44'h52621526856;
assign testcases[966] = 44'h63722107529;
assign testcases[967] = 44'h66312569512;
assign testcases[968] = 44'h63721625639;
assign testcases[969] = 44'h35122118934;
assign testcases[970] = 44'h82811108756;
assign testcases[971] = 44'h82811108756;
assign testcases[972] = 44'h83822107638;
assign testcases[973] = 44'h62712107a36;
assign testcases[974] = 44'h62752108739;
assign testcases[975] = 44'h43512848922;
assign testcases[976] = 44'h43512848922;
assign testcases[977] = 44'h55523769522;
assign testcases[978] = 44'h33531215727;
assign testcases[979] = 44'hb4812008535;
assign testcases[980] = 44'h64511219745;
assign testcases[981] = 44'h78412318634;
assign testcases[982] = 44'h44512b4585b;
assign testcases[983] = 44'h64511219745;
assign testcases[984] = 44'hb4812008535;
assign testcases[985] = 44'h45011107927;
assign testcases[986] = 44'h72611005627;
assign testcases[987] = 44'h43512848922;
assign testcases[988] = 44'h43212417522;
assign testcases[989] = 44'h72612316526;
assign testcases[990] = 44'h43212417522;
assign testcases[991] = 44'h42412748912;
assign testcases[992] = 44'h33212726812;
assign testcases[993] = 44'h42412748912;
assign testcases[994] = 44'h8372245b512;
assign testcases[995] = 44'h45112428834;
assign testcases[996] = 44'h16012004c3b;
assign testcases[997] = 44'h16012004c3b;
assign testcases[998] = 44'h68511106512;
assign testcases[999] = 44'h3601110292b;


  
  localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
  wire [$clog2(CLASS_CNT)-1:0] prediction;

  // Instantiate module under test
 winequality_red_ts #(
 ) dut (
    .data(data),
    .clk(clk),
    .rst(rst),
    .prediction(prediction)
  );
  
  always #halfT clk <= ~clk;

  integer i;
  initial begin
    $write("["); //" 
    for(i=0;i<TEST_CNT;i=i+1)
        runtestcase(i);
    $display("]");
    $finish;
  end

  task runtestcase(input integer i); begin
    data <= testcases[i];
    rst <= 1;
    clk <= 0;
    #period
    rst <= 0;
    #period
    #((FEAT_CNT+HIDDEN_CNT-1)*period)
    $write("%d, ",prediction);
  end
  endtask

endmodule
