












module cardio_bs #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 5


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 760'b1011011011110011000110010101010010110000110010001000101011100100100111011000001000000101010011011001001000101001011001011100110110001010111001000001110110010110001111100101110100100001011010001100100011011011101001001110000110110100100111010010000101000100000001000111011100110101110010011001101101011100110110111010010110001111111111100100010000111101100000110011001001010100000000111110000000001101010110001011001011000101101110011001010100011010000100000111000010100000111001101011001111010010001101000101000110011001010011001001001110110010100101000101001111111010010000100010001000010111101000001100000110000010101011100100100000110010101011011001100111100101100011111101001011011000100000011100110110001010100101100001011001110001010110101010100100011100 ;
  localparam Weights1 = 120'b110011011000011011101100100111001101001011100101100101101110110011011000110100111001110001000100110000001111100000010101 ;

  localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
  wire [SUM_BITS*CLASS_CNT-1:0] sums;

  seqlego #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) layers (
    .clk(clk),
    .rst(rst),
    .data(data),
    .out(sums)
  );

  argmax #(.SIZE(CLASS_CNT),.I($clog2(CLASS_CNT)),.K(SUM_BITS)) result (
     .inx(sums),
     .outimax(prediction)
  );

endmodule
