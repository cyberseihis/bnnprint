
















module winered_bnn1_bnnpaarter #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 4656'h0021002a00010021002a0000000d004e0001000d004a0001002600470001001d00460001001700450001002700440001000f004000010019003f0001001e003e0001002b003c00010024003b00010027003a0001002000380001001a00370001002100360001002500320001001e003100010018003000010017002e00010014002d00010014002c0001002500290001001400290001001f00230001001e002200010022003d0000001900330000001800310000001a003000000025002f00000014002f00000012002e0000001d002c0000002000290000001c00280000001000280000001c00240000001800240000001d00230000001400230000001b00220000001e00210000001a00200000001200200000000d001c00000014001a00000010001900000010001400000014002d0000001a002b0000001d00280000001000270000001f00230000001e00220000001a001d00000017001c0000001200260001001400170001001000170001001a001f00000019001c0000000f001b0000000d000f0000001700180000001800190001001200130001000f00130001000e00160000000c00110000000e001600010012001b0001001200140000001100160001000c00110001001100160000000d00100001000c000e0001000500150000000d00100000000500150001000d000f00010005000b0000000f001300000009000a0001000000080001000c000e00000001000400010002000700000003000600000005000b00010002000700010003000600010001000400000009000a0000000000080000 ;
localparam YMAP = 1280'h000000580001005d0000005500010051000100500001006a000100520001005c000000640000005f000100490001005600000062000100680000005e00010067000000610001005b000000540000006000000042000100390001005700000069000000530001004300000059000100340001004b0000006b000100410001005a0001006500010066000100350000004c00010063000100480001004f0001004d;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 240'b101011110101010111101111010101000101111001101110110011111110010011110100100011101000101011111101111001010101001011000101101011100011011000100010000100100000001111000110100000011011100000011101001111010010001011110000001101110000010000111001 ;
localparam WIDTH = 320'h07070707070607070706060706070707070707070707070707060707060707070706060707070707;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;
generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam subad = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(subad)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] < 0;
    initial begin
        #20
        $display("%b, %d | %d", signy, ymap, node[ymap]);
    end
end
endgenerate

initial begin
    #10
    for(j=0;j<FULLCNT;j=j+1) begin
        $display("%d | %d | %b, %d, %d", j, node[j], PAAR0[(j- FEAT_CNT )*48],  PAAR0[(j-FEAT_CNT)*48+16+:16], PAAR0[(j-FEAT_CNT)*48+32+:16]);
    end
end

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wneur[j])
            tmpscore = tmpscore + hidden[j];
        else 
            tmpscore = tmpscore + hidden_n[j];
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = tmpscore;
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
