module demox(input [111:0] a, output [15:0] o);
wire signed [10:0] t [15:0];
assign t[0] = + a[6:0] + a[13:7] - a[20:14] - a[27:21] - a[34:28] - a[41:35] - a[48:42] - a[55:49] - a[62:56] - a[69:63] + a[76:70] - a[83:77] - a[90:84] - a[97:91] - a[104:98] - a[111:105];assign o[0] = -220 < t[0];
assign t[1] = + a[6:0] + a[13:7] - a[20:14] - a[27:21] - a[34:28] - a[41:35] - a[48:42] + a[55:49] + a[62:56] - a[69:63] + a[76:70] + a[83:77] + a[90:84] + a[97:91] + a[104:98] - a[111:105];assign o[1] = 114 < t[1];
assign t[2] = - a[6:0] + a[13:7] - a[20:14] + a[27:21] + a[34:28] + a[41:35] - a[48:42] - a[55:49] + a[62:56] - a[69:63] + a[76:70] + a[83:77] - a[90:84] + a[97:91] - a[104:98] + a[111:105];assign o[2] = -45 < t[2];
assign t[3] = + a[6:0] - a[13:7] - a[20:14] - a[27:21] + a[34:28] - a[41:35] + a[48:42] + a[55:49] + a[62:56] + a[69:63] + a[76:70] - a[83:77] + a[90:84] + a[97:91] - a[104:98] + a[111:105];assign o[3] = 196 < t[3];
assign t[4] = + a[6:0] - a[13:7] + a[20:14] - a[27:21] - a[34:28] + a[41:35] - a[48:42] + a[55:49] - a[62:56] - a[69:63] + a[76:70] + a[83:77] - a[90:84] + a[97:91] - a[104:98] + a[111:105];assign o[4] = -183 < t[4];
assign t[5] = - a[6:0] + a[13:7] - a[20:14] + a[27:21] + a[34:28] + a[41:35] + a[48:42] - a[55:49] + a[62:56] - a[69:63] + a[76:70] + a[83:77] - a[90:84] + a[97:91] + a[104:98] + a[111:105];assign o[5] = 299 < t[5];
assign t[6] = + a[6:0] + a[13:7] + a[20:14] + a[27:21] - a[34:28] + a[41:35] - a[48:42] + a[55:49] + a[62:56] + a[69:63] + a[76:70] + a[83:77] + a[90:84] - a[97:91] - a[104:98] - a[111:105];assign o[6] = 435 < t[6];
assign t[7] = + a[6:0] + a[13:7] + a[20:14] + a[27:21] + a[34:28] + a[41:35] - a[48:42] - a[55:49] - a[62:56] - a[69:63] - a[76:70] - a[83:77] - a[90:84] + a[97:91] + a[104:98] + a[111:105];assign o[7] = 102 < t[7];
assign t[8] = + a[6:0] + a[13:7] - a[20:14] - a[27:21] - a[34:28] - a[41:35] - a[48:42] - a[55:49] - a[62:56] + a[69:63] - a[76:70] + a[83:77] - a[90:84] - a[97:91] + a[104:98] - a[111:105];assign o[8] = -267 < t[8];
assign t[9] = + a[6:0] - a[13:7] + a[20:14] - a[27:21] + a[34:28] + a[41:35] + a[48:42] + a[55:49] - a[62:56] + a[69:63] + a[76:70] + a[83:77] - a[90:84] + a[97:91] + a[104:98] + a[111:105];assign o[9] = 236 < t[9];
assign t[10] = - a[6:0] + a[13:7] - a[20:14] - a[27:21] - a[34:28] + a[41:35] + a[48:42] + a[55:49] - a[62:56] + a[69:63] - a[76:70] + a[83:77] - a[90:84] - a[97:91] + a[104:98] - a[111:105];assign o[10] = -75 < t[10];
assign t[11] = - a[6:0] - a[13:7] - a[20:14] + a[27:21] + a[34:28] + a[41:35] + a[48:42] + a[55:49] - a[62:56] - a[69:63] - a[76:70] - a[83:77] - a[90:84] - a[97:91] + a[104:98] - a[111:105];assign o[11] = 91 < t[11];
assign t[12] = - a[6:0] + a[13:7] + a[20:14] - a[27:21] - a[34:28] + a[41:35] + a[48:42] + a[55:49] + a[62:56] - a[69:63] + a[76:70] + a[83:77] - a[90:84] + a[97:91] + a[104:98] - a[111:105];assign o[12] = 203 < t[12];
assign t[13] = + a[6:0] + a[13:7] - a[20:14] - a[27:21] - a[34:28] - a[41:35] - a[48:42] - a[55:49] + a[62:56] + a[69:63] - a[76:70] + a[83:77] + a[90:84] + a[97:91] + a[104:98] + a[111:105];assign o[13] = 154 < t[13];
assign t[14] = + a[6:0] - a[13:7] + a[20:14] - a[27:21] - a[34:28] + a[41:35] + a[48:42] + a[55:49] + a[62:56] + a[69:63] - a[76:70] + a[83:77] + a[90:84] - a[97:91] + a[104:98] - a[111:105];assign o[14] = 22 < t[14];
assign t[15] = + a[6:0] + a[13:7] + a[20:14] + a[27:21] + a[34:28] + a[41:35] + a[48:42] + a[55:49] + a[62:56] + a[69:63] + a[76:70] - a[83:77] + a[90:84] - a[97:91] - a[104:98] - a[111:105];assign o[15] = 646 < t[15];
endmodule
