`timescale 1us/1ns









module tbpendigits_tnn1_tnnpar #(

parameter FEAT_CNT = 16,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 10,
parameter TEST_CNT = 1000


)();
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
reg clk;
reg [FEAT_CNT*FEAT_BITS-1:0] features;
wire [$clog2(CLASS_CNT)-1:0] prediction;
wire [FEAT_CNT*FEAT_BITS-1:0] testcases [TEST_CNT-1:0];
parameter Nsperiod=5000;
localparam period=Nsperiod/500;


assign testcases[0] = 64'hf6ef89400469d4f8;
assign testcases[1] = 64'h1f0b062275c7f4e0;
assign testcases[2] = 64'h034488ccffecb590;
assign testcases[3] = 64'h0b4c7f5e73b1f1f0;
assign testcases[4] = 64'h083566aaddffd8b0;
assign testcases[5] = 64'h333c063083c8feff;
assign testcases[6] = 64'h0b8afcbf6e64c0f0;
assign testcases[7] = 64'h90f6fe7f0a12a060;
assign testcases[8] = 64'hfff5a031096c82e2;
assign testcases[9] = 64'he4ec8f2c0450c4f9;
assign testcases[10] = 64'h030d6fdfaab0f5ec;
assign testcases[11] = 64'he0ffbd53034eaaf8;
assign testcases[12] = 64'h00032a8d95c6fcff;
assign testcases[13] = 64'h031d6fbd94e0f9cf;
assign testcases[14] = 64'h4f48092d8eedf6e0;
assign testcases[15] = 64'h30051d6dbbfff9c6;
assign testcases[16] = 64'h10082f7f88ccfbd8;
assign testcases[17] = 64'h30094fafbdc4fadf;
assign testcases[18] = 64'h0f09230045a9f7b4;
assign testcases[19] = 64'h0f073185cbfcf3c0;
assign testcases[20] = 64'hfff4a030086ca3c2;
assign testcases[21] = 64'h0e4c8ecfffeca870;
assign testcases[22] = 64'hfff5b041055bb5e2;
assign testcases[23] = 64'hfe98220f6dc0f8ac;
assign testcases[24] = 64'h36774f0b2071c5f9;
assign testcases[25] = 64'h0b5bbcaf8e72b0f2;
assign testcases[26] = 64'hf6ed7f1c0460d1f6;
assign testcases[27] = 64'h004498dbcfa5d2f7;
assign testcases[28] = 64'hbf75110d77d0f99a;
assign testcases[29] = 64'h00306282b1e0f5df;
assign testcases[30] = 64'ha0993f087dfff895;
assign testcases[31] = 64'hfff7c140064db8f6;
assign testcases[32] = 64'h5f6844097bedf6f0;
assign testcases[33] = 64'hc0f7df6f0b0370c4;
assign testcases[34] = 64'hadd9fddf8e5a2500;
assign testcases[35] = 64'h10093f6c88ccfbe5;
assign testcases[36] = 64'hfff6c030056b92f5;
assign testcases[37] = 64'h087caf5d5190f6fc;
assign testcases[38] = 64'h046fbfb2febfb0fa;
assign testcases[39] = 64'h0f08105389def8f1;
assign testcases[40] = 64'h6e6206187bcffaf0;
assign testcases[41] = 64'hfff7a230087b93e5;
assign testcases[42] = 64'h22695f0b0260c3fa;
assign testcases[43] = 64'h02082f7cbafef5d0;
assign testcases[44] = 64'h00265a9cdffef7e1;
assign testcases[45] = 64'h916c1f0450b4fbff;
assign testcases[46] = 64'h20061d4f8bcefce8;
assign testcases[47] = 64'h0f1810247accf7c5;
assign testcases[48] = 64'hfff4b142065990e0;
assign testcases[49] = 64'h004589cdcfabc6fa;
assign testcases[50] = 64'h00092f6e98ddf9f2;
assign testcases[51] = 64'h003265a9ddfffbc8;
assign testcases[52] = 64'hc3f9bf4e0640c3f9;
assign testcases[53] = 64'h033668acdfffe8c0;
assign testcases[54] = 64'h0c8bfcaf6c61c0f3;
assign testcases[55] = 64'hfff8e0500568c3f7;
assign testcases[56] = 64'h20073e8d9bdffad3;
assign testcases[57] = 64'h0f18302278ccf6c2;
assign testcases[58] = 64'hd1f8bf4f0942c0c3;
assign testcases[59] = 64'h21684f084091e7ff;
assign testcases[60] = 64'hbf61003f86f0ffa9;
assign testcases[61] = 64'h00095f97e6fffed5;
assign testcases[62] = 64'h80f2fbaf4f0730a2;
assign testcases[63] = 64'h000a4f7886dcf8d0;
assign testcases[64] = 64'h78510256aafffaf0;
assign testcases[65] = 64'h9f66100867c4fbdf;
assign testcases[66] = 64'h00076c95e8fffdf6;
assign testcases[67] = 64'h60783d074395d9ff;
assign testcases[68] = 64'hdf87300b59a2f6df;
assign testcases[69] = 64'hd0fdcf74042f9cd0;
assign testcases[70] = 64'h10082f8ddad9f6fd;
assign testcases[71] = 64'hb1f8ef7f1a0270c6;
assign testcases[72] = 64'h0b7c7f5f5760c3f5;
assign testcases[73] = 64'h094b9ddfffdbc5c0;
assign testcases[74] = 64'h003a8fad82e4ffbe;
assign testcases[75] = 64'h7f76430568bbf7f0;
assign testcases[76] = 64'hf5fcaf3d0730a1f6;
assign testcases[77] = 64'h12593f083090e6fc;
assign testcases[78] = 64'h00082f7e99effbd4;
assign testcases[79] = 64'h20072f7fbbfff8c1;
assign testcases[80] = 64'h0f0a25002589f9c5;
assign testcases[81] = 64'h094c8f7b74a0e3f7;
assign testcases[82] = 64'h2f18200769dcfcb7;
assign testcases[83] = 64'h033a1f063080c2f5;
assign testcases[84] = 64'hfff8d0610468a1e3;
assign testcases[85] = 64'hffd271023e9e90e3;
assign testcases[86] = 64'h675f0c3a8beff9f0;
assign testcases[87] = 64'ha1f7df5f0830b0f8;
assign testcases[88] = 64'hd3fabf4e0730b186;
assign testcases[89] = 64'h00469befecc3f8ff;
assign testcases[90] = 64'hfff7b350004690e3;
assign testcases[91] = 64'h917b3f083080d4f6;
assign testcases[92] = 64'h0b5cad6f5850b0f4;
assign testcases[93] = 64'h70785f0c4dbdf8f0;
assign testcases[94] = 64'h0f3d7dacecfad6a0;
assign testcases[95] = 64'hf5fcbf5e090270d3;
assign testcases[96] = 64'h09497abdfffdd6a0;
assign testcases[97] = 64'h0f8f9ac0fbbf83c6;
assign testcases[98] = 64'h344c0a014084caff;
assign testcases[99] = 64'h0f060048affce395;
assign testcases[100] = 64'hd0f7de6f0c2481f2;
assign testcases[101] = 64'h00083f8f87cbfae3;
assign testcases[102] = 64'hc1f9af3f0a43b0f1;
assign testcases[103] = 64'hf3ff9c50022e8ad7;
assign testcases[104] = 64'ha0f4fcaf2f0822a1;
assign testcases[105] = 64'h00092f5b99dffef6;
assign testcases[106] = 64'hb5fbbf4e0730a294;
assign testcases[107] = 64'h83f8ff6f0a1290f4;
assign testcases[108] = 64'hfff7d0610368b2f7;
assign testcases[109] = 64'h0e4d9f8e71b3f6e0;
assign testcases[110] = 64'h01757f1b2090f6fc;
assign testcases[111] = 64'hb3f7ce6f0d0550c2;
assign testcases[112] = 64'h608b3f084091d5fe;
assign testcases[113] = 64'he1ffbd55075cb4e0;
assign testcases[114] = 64'h001b8ecfe7ffbcf8;
assign testcases[115] = 64'h03578e7f5870d1f7;
assign testcases[116] = 64'hfff7a121066890f1;
assign testcases[117] = 64'h454c062083c8ffcf;
assign testcases[118] = 64'h1f18000148adfbb7;
assign testcases[119] = 64'h40084fbdf4fc98f6;
assign testcases[120] = 64'hc0fd88100d6ad6ef;
assign testcases[121] = 64'hfff472035ebca0f7;
assign testcases[122] = 64'ha0f6df5f0931b2f7;
assign testcases[123] = 64'hc0f5ed9f3e0752b2;
assign testcases[124] = 64'he1fabf4f083091d8;
assign testcases[125] = 64'h0e4f8f6f5791c0f3;
assign testcases[126] = 64'h054497dbfff8f0f4;
assign testcases[127] = 64'h20072e7f79befcf8;
assign testcases[128] = 64'h00469befffc8f8ff;
assign testcases[129] = 64'h0f18102267bbf9c5;
assign testcases[130] = 64'hfff8c0420667a1f2;
assign testcases[131] = 64'h000bafb9fbaf85e8;
assign testcases[132] = 64'he9bf5f0a0270d4fb;
assign testcases[133] = 64'h5047071172c5faff;
assign testcases[134] = 64'hd7bf3f0840c2f9bf;
assign testcases[135] = 64'h414f0f2370c3f9fd;
assign testcases[136] = 64'h405a1f064294d8ff;
assign testcases[137] = 64'h086abdfffec99570;
assign testcases[138] = 64'h065bbf8f6790e5fb;
assign testcases[139] = 64'h46cdfd9f1800a5ec;
assign testcases[140] = 64'h81f4fb9f1d0560d4;
assign testcases[141] = 64'h616c3f074082d8fe;
assign testcases[142] = 64'h0f0a103077ccfad6;
assign testcases[143] = 64'h00367bbfebd3fbef;
assign testcases[144] = 64'hfff4b0520748a3f5;
assign testcases[145] = 64'h40070f6fccfff7c0;
assign testcases[146] = 64'h074a9defffda9570;
assign testcases[147] = 64'h0c4e8f8f6780c1f3;
assign testcases[148] = 64'h2f2b150052b4f3b0;
assign testcases[149] = 64'h0f6f5f383083d6f8;
assign testcases[150] = 64'h004488ccffdfaa65;
assign testcases[151] = 64'h0d4b8ccefffdc7a0;
assign testcases[152] = 64'h1f13032d9fffd880;
assign testcases[153] = 64'h70894f0a2180d4fa;
assign testcases[154] = 64'h004175baffffd2de;
assign testcases[155] = 64'h086ccdb0f4ffb8d2;
assign testcases[156] = 64'hf1fca844085f98d0;
assign testcases[157] = 64'h0d4f5e4660a2d6fc;
assign testcases[158] = 64'h7f75510569cefbf0;
assign testcases[159] = 64'h00081f6ea9effbd6;
assign testcases[160] = 64'h042a5d8fafdffcf0;
assign testcases[161] = 64'h0367bdb1f3ffcc90;
assign testcases[162] = 64'h705b1f086accf5e0;
assign testcases[163] = 64'h0f5fbfcf9f84c0f2;
assign testcases[164] = 64'h20082f7fabfef6c3;
assign testcases[165] = 64'hf7ce5f0b0460d2f8;
assign testcases[166] = 64'h6c5003368acffff4;
assign testcases[167] = 64'h003888a1e8ffffe7;
assign testcases[168] = 64'hf1ff89110b79e0f9;
assign testcases[169] = 64'h20082f6e9cdffed7;
assign testcases[170] = 64'h12655f0830a2f7fd;
assign testcases[171] = 64'hffe7a040033a83c4;
assign testcases[172] = 64'h0f150056a9fdeca6;
assign testcases[173] = 64'hfff7b120068890f2;
assign testcases[174] = 64'h014488cbffffc7a0;
assign testcases[175] = 64'h0f2f6d9bcafae8b0;
assign testcases[176] = 64'h0f4f8ecefefad3b0;
assign testcases[177] = 64'h00196fbffeccd7fe;
assign testcases[178] = 64'h0b5daf5d4480d3f5;
assign testcases[179] = 64'hfff69001098c92f4;
assign testcases[180] = 64'h08589bdefff9f3c0;
assign testcases[181] = 64'h888f4f0e6fdef7f0;
assign testcases[182] = 64'h7f7440085bbefef3;
assign testcases[183] = 64'hf6ed8f3c0540a1f5;
assign testcases[184] = 64'h00174c8ecffff9c3;
assign testcases[185] = 64'h445f1f044083c8ff;
assign testcases[186] = 64'h00367ccffbf2b3cd;
assign testcases[187] = 64'h303909004094d9ff;
assign testcases[188] = 64'h044b8fcaf0ffc6e3;
assign testcases[189] = 64'hb1f6fe9f2c055093;
assign testcases[190] = 64'h0c5caeffb9c0f7ed;
assign testcases[191] = 64'h5f59610437a9f7f0;
assign testcases[192] = 64'h0b4d7fbfeffedab0;
assign testcases[193] = 64'hfadf7f2b0540b1f5;
assign testcases[194] = 64'h00073d8f98d7fbff;
assign testcases[195] = 64'he8cf5f1b0350b3f8;
assign testcases[196] = 64'h00074c9ca6e4faff;
assign testcases[197] = 64'h1f003b8cdeffb985;
assign testcases[198] = 64'h100a5fcfcdc3f6ee;
assign testcases[199] = 64'h094c8f6b61a0d6fb;
assign testcases[200] = 64'h0377ebdfbc90c4f8;
assign testcases[201] = 64'h0557a9fd9f96c0f4;
assign testcases[202] = 64'hfff8c170012986d0;
assign testcases[203] = 64'h0f0710478ccffff8;
assign testcases[204] = 64'h4048062072b6fbff;
assign testcases[205] = 64'hf4de6a0a3f87e0f9;
assign testcases[206] = 64'h1f092578ccf9e4a0;
assign testcases[207] = 64'h09398bcdfffbd5c0;
assign testcases[208] = 64'h0a4c9edfffdaa480;
assign testcases[209] = 64'h00083f7f88cefee6;
assign testcases[210] = 64'hd0fbb952084fbaec;
assign testcases[211] = 64'h00459adfae96c5fb;
assign testcases[212] = 64'h6f5523087cdff9e0;
assign testcases[213] = 64'h0021457999bcefff;
assign testcases[214] = 64'hfff8f061034aa6f8;
assign testcases[215] = 64'h053677aaddfff7f0;
assign testcases[216] = 64'hfff6b051055ba5c2;
assign testcases[217] = 64'hf4ff99400784f3fd;
assign testcases[218] = 64'hfff8c3500236a3d6;
assign testcases[219] = 64'h0e5e9f6b7380c5f8;
assign testcases[220] = 64'h00564f083193f6fc;
assign testcases[221] = 64'h0f072267aceef8e0;
assign testcases[222] = 64'h00082f6f9ceffdd7;
assign testcases[223] = 64'h0f4f5f274084cafd;
assign testcases[224] = 64'h0e6bdebfaf91e0f8;
assign testcases[225] = 64'hdf85200b6ac3fcbf;
assign testcases[226] = 64'h807b3f084295ebff;
assign testcases[227] = 64'h1f0a34003699f8a5;
assign testcases[228] = 64'hfff6a1100477c2f6;
assign testcases[229] = 64'hfff8e250034984f4;
assign testcases[230] = 64'h40592f073183d8ff;
assign testcases[231] = 64'h7f79630749baf6f0;
assign testcases[232] = 64'h6f58500557c8f4d0;
assign testcases[233] = 64'h05488acdffeab580;
assign testcases[234] = 64'h6b530759acfff8f0;
assign testcases[235] = 64'h00182f39a9f9a692;
assign testcases[236] = 64'h10062c6faccdfdf7;
assign testcases[237] = 64'hf9efa751065ab6b0;
assign testcases[238] = 64'h034a8fdff8e0a5cf;
assign testcases[239] = 64'hd0f8cf5f0a0170c5;
assign testcases[240] = 64'h30072e8f89cffdd8;
assign testcases[241] = 64'hf8ff9f3c063091f5;
assign testcases[242] = 64'h6f78440669ccf7f0;
assign testcases[243] = 64'haf57001b76d4ffcf;
assign testcases[244] = 64'h0f38411047c9f4a1;
assign testcases[245] = 64'h001a7fabf6ffbdfa;
assign testcases[246] = 64'h128cdf5e0270e8fc;
assign testcases[247] = 64'h8cc7faefaf5b2600;
assign testcases[248] = 64'h0e5faea2d0facf98;
assign testcases[249] = 64'h05478ccfffd8a070;
assign testcases[250] = 64'h095aae7f7470b7fc;
assign testcases[251] = 64'h80893d0540a5fbff;
assign testcases[252] = 64'h100a4f7987ddf6d0;
assign testcases[253] = 64'h0f090449adfbf4c0;
assign testcases[254] = 64'h303708025296cbff;
assign testcases[255] = 64'h73f5ed6f0931c0f4;
assign testcases[256] = 64'h760660a6fd9ce2ff;
assign testcases[257] = 64'hc2f9cf5d0550c3fb;
assign testcases[258] = 64'hf8bd61054f95f0fe;
assign testcases[259] = 64'h00468ceff9d0c5dc;
assign testcases[260] = 64'h20072f8f88cdfbd5;
assign testcases[261] = 64'hd1fecf66031f7cb0;
assign testcases[262] = 64'h6046043283c6faff;
assign testcases[263] = 64'h40675f0f1967c9fe;
assign testcases[264] = 64'h3f1800458bdff9c4;
assign testcases[265] = 64'hf0f9bf5f091181e5;
assign testcases[266] = 64'h0f5f9c90e1fbcf7a;
assign testcases[267] = 64'h0a498bcdfffef7e0;
assign testcases[268] = 64'ha3f8df5f0820a1c6;
assign testcases[269] = 64'hc0fccf64044ea4d9;
assign testcases[270] = 64'hffa5410b5da3f0ec;
assign testcases[271] = 64'h0e4f7f4a5290d1f0;
assign testcases[272] = 64'h0e6f7f584062b7fb;
assign testcases[273] = 64'h01483f0a3290f4fa;
assign testcases[274] = 64'h455d1d0450b3f8ff;
assign testcases[275] = 64'h0b4d8f6971b0f1f2;
assign testcases[276] = 64'ha0f5ed7f0c0480f2;
assign testcases[277] = 64'h04002679bcffca94;
assign testcases[278] = 64'h0f1800378bfdf8d7;
assign testcases[279] = 64'h3f37061c7ddcf5d0;
assign testcases[280] = 64'h40073f7dbffef4d5;
assign testcases[281] = 64'h0e8dfc8f4b40b0f7;
assign testcases[282] = 64'h20063b8ceeeafbff;
assign testcases[283] = 64'h30472d074496daff;
assign testcases[284] = 64'h10064b8883d4f9ff;
assign testcases[285] = 64'h3f09313087eaf5b6;
assign testcases[286] = 64'h415b1d034084c9ff;
assign testcases[287] = 64'h6d50071b7ddff8f0;
assign testcases[288] = 64'h204b1f035295eaff;
assign testcases[289] = 64'h10093f8c64d2f6ff;
assign testcases[290] = 64'h10083d8abdfff8c4;
assign testcases[291] = 64'h1f08003288dcf7b4;
assign testcases[292] = 64'h10073e8b72c3faff;
assign testcases[293] = 64'h845b0b1360b3e9ff;
assign testcases[294] = 64'h06489ccf8980c5fc;
assign testcases[295] = 64'h00083f7f8bcffcd6;
assign testcases[296] = 64'hc0a93c057beffa87;
assign testcases[297] = 64'h0f2a34357aebf5d0;
assign testcases[298] = 64'hfff79220086c94e5;
assign testcases[299] = 64'h20073e8cbdfff8d2;
assign testcases[300] = 64'h00085aa4e8ffffe9;
assign testcases[301] = 64'h6c530358adfff7f0;
assign testcases[302] = 64'h0a4d7f6a6390d3f8;
assign testcases[303] = 64'h30082f8c9beff7c2;
assign testcases[304] = 64'h00074c9cb6d4f9ff;
assign testcases[305] = 64'h0d4d8eceffca9550;
assign testcases[306] = 64'h0d16599edffcf4c0;
assign testcases[307] = 64'h00064a9994e5fbff;
assign testcases[308] = 64'hdf79071e78d0f8af;
assign testcases[309] = 64'h40094f96f1fdaa51;
assign testcases[310] = 64'h0e6f9f6a7070c5f7;
assign testcases[311] = 64'hc4661f076bcff6c0;
assign testcases[312] = 64'h20083f8ab6fcfff7;
assign testcases[313] = 64'h0e4c9decf6c0a7cf;
assign testcases[314] = 64'h10072d7faaeffbc5;
assign testcases[315] = 64'h35c4faaf1d0570e2;
assign testcases[316] = 64'h0f183276abfcf5e0;
assign testcases[317] = 64'h7f7741055abcf6d0;
assign testcases[318] = 64'h1f100666e4f992d3;
assign testcases[319] = 64'h0f120148a8f8f7a0;
assign testcases[320] = 64'h08388bcdffd8b0a6;
assign testcases[321] = 64'h0b5d9f6b60a0f4f2;
assign testcases[322] = 64'h7f7826086adcf7e0;
assign testcases[323] = 64'h59340a5daffef7e0;
assign testcases[324] = 64'he0fbbf58065bb4c9;
assign testcases[325] = 64'h044688ccfffcc680;
assign testcases[326] = 64'h00094fbef9b7f3f7;
assign testcases[327] = 64'hc0f7df5f0a1290f4;
assign testcases[328] = 64'h825c0c0260b4fbff;
assign testcases[329] = 64'h14674f0740a3f9c6;
assign testcases[330] = 64'hfcca50055eb5efb4;
assign testcases[331] = 64'h0f1b35303488f9f6;
assign testcases[332] = 64'h00094f7e89cdf8e1;
assign testcases[333] = 64'hcf8620095ea7f1ff;
assign testcases[334] = 64'h0f2a3471a7eaf4e0;
assign testcases[335] = 64'hfff381004accb1f7;
assign testcases[336] = 64'h10093f6988cffad4;
assign testcases[337] = 64'h03574f0740a1f7ff;
assign testcases[338] = 64'h12092f7faaedf6d0;
assign testcases[339] = 64'h0f081156aafaf4c0;
assign testcases[340] = 64'h0f0914478ac9f6f0;
assign testcases[341] = 64'h304a1e054284c9ff;
assign testcases[342] = 64'h1f1b050052b4f3d1;
assign testcases[343] = 64'hfabf6f1b0340a3e8;
assign testcases[344] = 64'hbf67000b4aa3f8de;
assign testcases[345] = 64'h50095fdfe4fcb8f6;
assign testcases[346] = 64'h7f65220558bbfaf0;
assign testcases[347] = 64'hfff59322086b92b0;
assign testcases[348] = 64'h086ace9f7960a8fc;
assign testcases[349] = 64'h00194f8fa8defad6;
assign testcases[350] = 64'h0a29699bddffe7c0;
assign testcases[351] = 64'h0f4c8ccdfff8c0a7;
assign testcases[352] = 64'h40481c054397dcff;
assign testcases[353] = 64'h002a8fefcea5f9ff;
assign testcases[354] = 64'h71d5fcbf4e082190;
assign testcases[355] = 64'h0c0310488ddffae3;
assign testcases[356] = 64'hd0f6dc7f1d063082;
assign testcases[357] = 64'h0f3950316bcffbc5;
assign testcases[358] = 64'hef98500063c2f8ce;
assign testcases[359] = 64'h61f5fd7f0a01a0e4;
assign testcases[360] = 64'h0f18102057baf6b2;
assign testcases[361] = 64'h213b0c034093e8ff;
assign testcases[362] = 64'h445e1f063081d5fd;
assign testcases[363] = 64'h0b5abdfffdd7b190;
assign testcases[364] = 64'h8f87430468ccf8d0;
assign testcases[365] = 64'h0e6fcfcbb0f1fcbf;
assign testcases[366] = 64'h0f29223065bafac6;
assign testcases[367] = 64'h0f18100149bcf7c4;
assign testcases[368] = 64'h0c5c7f3c3360b1f2;
assign testcases[369] = 64'hfff7c032088ab2f3;
assign testcases[370] = 64'h00082f6ebaeff9d3;
assign testcases[371] = 64'h0a69dafaaf94d0f6;
assign testcases[372] = 64'h0f09024487d8f4d0;
assign testcases[373] = 64'h1f08311056abfbd5;
assign testcases[374] = 64'hfea6400557b0f4ff;
assign testcases[375] = 64'hfff6b220068a71e3;
assign testcases[376] = 64'h84f7fe8f0c0470f3;
assign testcases[377] = 64'hfebf670b5da3f0fc;
assign testcases[378] = 64'h30084f9e97def8c3;
assign testcases[379] = 64'hb0f6dd6f0c2480e1;
assign testcases[380] = 64'h5f55300759adfbf0;
assign testcases[381] = 64'h10061c5f9bcdfcf6;
assign testcases[382] = 64'h435d2f073180c2f5;
assign testcases[383] = 64'h9b7100258bfff6c2;
assign testcases[384] = 64'h0f09120046aafcc9;
assign testcases[385] = 64'h0b4b8dcfffcb9660;
assign testcases[386] = 64'h0368cd9f87a0e9fe;
assign testcases[387] = 64'hc1f8cf5f0a32a0e1;
assign testcases[388] = 64'h06487cafeff9f1f0;
assign testcases[389] = 64'h454b2b0599fff8f0;
assign testcases[390] = 64'h11483f073080c3f8;
assign testcases[391] = 64'he5de6f0b2290f5ca;
assign testcases[392] = 64'h030c3f7bb8f9f2d0;
assign testcases[393] = 64'hcc99400a5cc4f9bf;
assign testcases[394] = 64'h40591c044093e9ff;
assign testcases[395] = 64'h4339062071b5eaff;
assign testcases[396] = 64'hf5fcaf4f081280d4;
assign testcases[397] = 64'hd0fcbf68020d6cc6;
assign testcases[398] = 64'h0f4950326abffcd6;
assign testcases[399] = 64'h10093f7d88dcf8c4;
assign testcases[400] = 64'h100a4f7da9effae2;
assign testcases[401] = 64'h095aadffeec1f0fd;
assign testcases[402] = 64'hfff8b343085892e0;
assign testcases[403] = 64'h024488ccfffcd6b0;
assign testcases[404] = 64'hf7ef6f0a0070d6fe;
assign testcases[405] = 64'h001a7fefc6f2fcaa;
assign testcases[406] = 64'h536c2f083081c5fc;
assign testcases[407] = 64'h10161f0c59c9f9a6;
assign testcases[408] = 64'h345e1f064091d6fd;
assign testcases[409] = 64'h00083f7f89cffbd7;
assign testcases[410] = 64'h6f6605299efff8f0;
assign testcases[411] = 64'hfcaf54003d9af8dc;
assign testcases[412] = 64'h0f084d8ccbfcfac0;
assign testcases[413] = 64'h0f08102479daf5a4;
assign testcases[414] = 64'h051e6b93e0f4fddf;
assign testcases[415] = 64'h002d9fabe5ffaec4;
assign testcases[416] = 64'h0f293300369af8c5;
assign testcases[417] = 64'h00185c98cffff8c2;
assign testcases[418] = 64'h094b9e7f4a71c0f1;
assign testcases[419] = 64'h09386aacdffff7f0;
assign testcases[420] = 64'h7f78430468dbf6f0;
assign testcases[421] = 64'hc0fbaf53056bc2f5;
assign testcases[422] = 64'h0b4d8f4b4081c4f9;
assign testcases[423] = 64'h10082f7e89ddf7d2;
assign testcases[424] = 64'h0167bf90d0ffcfc5;
assign testcases[425] = 64'h7f78240579ecf6f0;
assign testcases[426] = 64'hfcce66000f6fc5fa;
assign testcases[427] = 64'h00084c8681e2f8ff;
assign testcases[428] = 64'hf8fdaf3d081370e1;
assign testcases[429] = 64'h40061e6dbdfff8e8;
assign testcases[430] = 64'h53c3fbaf2e0650c1;
assign testcases[431] = 64'h9f55001682e2fcac;
assign testcases[432] = 64'h0e5daf7f6680d3f6;
assign testcases[433] = 64'h8d6407399cfff8f0;
assign testcases[434] = 64'h40885f0f0766caff;
assign testcases[435] = 64'hffd772002964b0f5;
assign testcases[436] = 64'h0f08114185d6f0d1;
assign testcases[437] = 64'h0a386cafeffbf5d0;
assign testcases[438] = 64'h0a7bec9f5e50a6f8;
assign testcases[439] = 64'hf6de5f0a31b0f6dd;
assign testcases[440] = 64'h10072d6facddfae4;
assign testcases[441] = 64'hd0f8cf5f0a2291e5;
assign testcases[442] = 64'h5f57320668c9f4d0;
assign testcases[443] = 64'h20072e6fabdcfbd7;
assign testcases[444] = 64'h00174e8faaedf9e2;
assign testcases[445] = 64'h0f7eddff9f75c0f2;
assign testcases[446] = 64'h00084e79c8feffe9;
assign testcases[447] = 64'h021c5c71b0f9fff5;
assign testcases[448] = 64'h474e0e2f8fddf7f0;
assign testcases[449] = 64'h7c54082b8eeff8f0;
assign testcases[450] = 64'h0f4e9f7b64a1f3f0;
assign testcases[451] = 64'h20043988d8fdfffb;
assign testcases[452] = 64'hf3facf4d0720a1f7;
assign testcases[453] = 64'h00368bdffdd6f6fc;
assign testcases[454] = 64'h08296baeeffdd6a0;
assign testcases[455] = 64'h033c7ea4c0f7fff6;
assign testcases[456] = 64'h1f08101369bcf9c5;
assign testcases[457] = 64'h425b1c014096ddff;
assign testcases[458] = 64'h20081f6ca8eef8c2;
assign testcases[459] = 64'h0a3768aadfffd8a0;
assign testcases[460] = 64'h0f28201157bbfef8;
assign testcases[461] = 64'h002679b4e9fffcd7;
assign testcases[462] = 64'h00297dbdffcae5fd;
assign testcases[463] = 64'h00266bbfefc9fcdf;
assign testcases[464] = 64'hd0660c178cfff8c5;
assign testcases[465] = 64'hbf78300769c5fcbe;
assign testcases[466] = 64'h0256bb8f6b60b1f5;
assign testcases[467] = 64'h695f2d087aecf5e0;
assign testcases[468] = 64'h6058081173c8feff;
assign testcases[469] = 64'h00082f8fcde6fcbf;
assign testcases[470] = 64'h0081e6fdaf2d0776;
assign testcases[471] = 64'h10483f093383c5fa;
assign testcases[472] = 64'h065caffdf4a099df;
assign testcases[473] = 64'h064eaffdf4a077af;
assign testcases[474] = 64'h7f61240a6fdff5e0;
assign testcases[475] = 64'h416d3f052074c9ff;
assign testcases[476] = 64'he89f2f0640b3f9cf;
assign testcases[477] = 64'h0f1800147afdf6d7;
assign testcases[478] = 64'h40d2fc7f0a11a0f4;
assign testcases[479] = 64'h0f0800358beff9b6;
assign testcases[480] = 64'h20095c95d6ffffe7;
assign testcases[481] = 64'h4239043072b6fbff;
assign testcases[482] = 64'h4f40071a8ceff8f0;
assign testcases[483] = 64'h20573f0a3283d8ff;
assign testcases[484] = 64'hfef0a0420c5fa9f1;
assign testcases[485] = 64'hf2fbbf5f082080e4;
assign testcases[486] = 64'hf7ed8f2e0843a0e3;
assign testcases[487] = 64'ha4f8fe9f3d063092;
assign testcases[488] = 64'h0e5f9c81d0f8ce7b;
assign testcases[489] = 64'hfff7a330087ab5f5;
assign testcases[490] = 64'h5d70310469cffff7;
assign testcases[491] = 64'h0c7dfeaf6c60c8ff;
assign testcases[492] = 64'h00094f9cbafef5c4;
assign testcases[493] = 64'h0f19125194f6f1c0;
assign testcases[494] = 64'h0f050248a9fad690;
assign testcases[495] = 64'h0b497bacefffd8a0;
assign testcases[496] = 64'hfff480041d9d81e0;
assign testcases[497] = 64'h0f051158acfbf1c0;
assign testcases[498] = 64'h01295c99cefff7e0;
assign testcases[499] = 64'hdaffbb65002497d8;
assign testcases[500] = 64'h00053aa8a3f5fbff;
assign testcases[501] = 64'h210d6fa5f4ed8820;
assign testcases[502] = 64'h5f57091b7deff8f0;
assign testcases[503] = 64'hd2fabf4e0730b0f7;
assign testcases[504] = 64'h6c5312086ddff9e0;
assign testcases[505] = 64'hfff692043ca990e2;
assign testcases[506] = 64'hfff370004baab1f5;
assign testcases[507] = 64'hd4fdbf7820096cb7;
assign testcases[508] = 64'h003276a9deffe5c5;
assign testcases[509] = 64'h076accff9f95d0f1;
assign testcases[510] = 64'h0e6f8f698082d8fb;
assign testcases[511] = 64'hcf78061f78c0f9bf;
assign testcases[512] = 64'h0f054379befff6e0;
assign testcases[513] = 64'h12074c87a0f1f9ff;
assign testcases[514] = 64'h8f77450b6eddf6d0;
assign testcases[515] = 64'h00003b7dcdfffec5;
assign testcases[516] = 64'h0c4d9ecf8a80d0f5;
assign testcases[517] = 64'h0f18211258caf6c0;
assign testcases[518] = 64'hf5df87200c6db3f2;
assign testcases[519] = 64'h004286cafeffc991;
assign testcases[520] = 64'h00180f1764c5f7c2;
assign testcases[521] = 64'hffd571012c8ac0e4;
assign testcases[522] = 64'h1f09021164d4f3a0;
assign testcases[523] = 64'h6f68520658baf8e0;
assign testcases[524] = 64'h0f00073eaeffed94;
assign testcases[525] = 64'hb9af3f0a1370d2f7;
assign testcases[526] = 64'h0f28101368bbf9c4;
assign testcases[527] = 64'hcf84100b75e2fca6;
assign testcases[528] = 64'h2f28200677f8c7d7;
assign testcases[529] = 64'hfff281001a9c80e3;
assign testcases[530] = 64'h4e4001167acffff1;
assign testcases[531] = 64'h0e5eaecf9d81d0f1;
assign testcases[532] = 64'hfff6a041045991d2;
assign testcases[533] = 64'h22695f0a0170c4fb;
assign testcases[534] = 64'h0f18203479ccf9d4;
assign testcases[535] = 64'h10082e6d9cdffdf8;
assign testcases[536] = 64'h6c600055aafff7f0;
assign testcases[537] = 64'hfece660646a0f6ff;
assign testcases[538] = 64'hc960011f7eb2f5bc;
assign testcases[539] = 64'hb8cf6f1b0450c0f6;
assign testcases[540] = 64'h0f3b7b9b6590c0f1;
assign testcases[541] = 64'hfff5a2022b9a90e3;
assign testcases[542] = 64'h6f6641096bcdf6c0;
assign testcases[543] = 64'h5f47061a7ddff9f0;
assign testcases[544] = 64'h03583f0740a1f5e9;
assign testcases[545] = 64'hf3eb9f3e0640b1f5;
assign testcases[546] = 64'h0f3b7d5f61a0d0f3;
assign testcases[547] = 64'hd8ff9f3b0270d5ed;
assign testcases[548] = 64'hf0ffaa510d6eb4e9;
assign testcases[549] = 64'h04477bafeff9f2f0;
assign testcases[550] = 64'h4f470a2d8feff7d0;
assign testcases[551] = 64'h0f5f7e4762b3f3f0;
assign testcases[552] = 64'h1f04387bcfffc890;
assign testcases[553] = 64'h0f3830559ceffbc7;
assign testcases[554] = 64'hffe8b062052b89d5;
assign testcases[555] = 64'h09295d8fafdffdf0;
assign testcases[556] = 64'h1f08004589ccf8f0;
assign testcases[557] = 64'h0f08103187f9f3a1;
assign testcases[558] = 64'h10071d9facfaff8d;
assign testcases[559] = 64'h0156adaf7980e3fa;
assign testcases[560] = 64'hffa7510849a3f0fc;
assign testcases[561] = 64'h10082f7f88dbf7c3;
assign testcases[562] = 64'h014a8fdce0fbcad4;
assign testcases[563] = 64'h0f0800278ceffac7;
assign testcases[564] = 64'hf6cf87300c5bb3f2;
assign testcases[565] = 64'hd0f7ee6f0c1592e6;
assign testcases[566] = 64'h00173e7bbefff9d7;
assign testcases[567] = 64'h00082f6e88cdf8e2;
assign testcases[568] = 64'h4249062062a5eaff;
assign testcases[569] = 64'h066acf8f74b0f8e8;
assign testcases[570] = 64'h094c8f7d5480c4f7;
assign testcases[571] = 64'h03546f2b3090f6ff;
assign testcases[572] = 64'he4ffbd570a5da6d0;
assign testcases[573] = 64'h10463d074295daff;
assign testcases[574] = 64'h0f0a032065b9f9f3;
assign testcases[575] = 64'hcf84200a68b1f8b9;
assign testcases[576] = 64'hfff78200077ab2f7;
assign testcases[577] = 64'h4f0b453057b9f6a5;
assign testcases[578] = 64'h0f2a432056baf6d1;
assign testcases[579] = 64'hffe472001a7da1f7;
assign testcases[580] = 64'h416b2f0640a3f8ff;
assign testcases[581] = 64'h30071f6f86cdfde5;
assign testcases[582] = 64'hc0f8ff9b44075b63;
assign testcases[583] = 64'hd0febd66063f9cc6;
assign testcases[584] = 64'hffaa51054fabe0fc;
assign testcases[585] = 64'h30082f9ffbd9f3fa;
assign testcases[586] = 64'h5f0f182057b8f4c4;
assign testcases[587] = 64'hc0f6fd9f2e0764e6;
assign testcases[588] = 64'hfcdf84041780f4ee;
assign testcases[589] = 64'h00093f8f99dffcca;
assign testcases[590] = 64'h00368aeec8c3faff;
assign testcases[591] = 64'hffa9440e6bb0f4ca;
assign testcases[592] = 64'h085baf7f74a0f5f4;
assign testcases[593] = 64'hffe590460d5da6d3;
assign testcases[594] = 64'h0d4c8ccefffec790;
assign testcases[595] = 64'hf7fe8f1c0460e1d6;
assign testcases[596] = 64'h0b4c8f9a80c0f6f3;
assign testcases[597] = 64'hb0f8ff6f0810b3c8;
assign testcases[598] = 64'h40062e8c74c3faef;
assign testcases[599] = 64'h10081f6f88dbf8d3;
assign testcases[600] = 64'h474f0c034082c5fb;
assign testcases[601] = 64'h0f5eaefdf5c0c8ee;
assign testcases[602] = 64'h0c6dbfaf9780c6fc;
assign testcases[603] = 64'h0f092367a9faf3d0;
assign testcases[604] = 64'hfaa640055ba6f6ff;
assign testcases[605] = 64'hf5ed7f0c0460d2e5;
assign testcases[606] = 64'hfff59232076a90e2;
assign testcases[607] = 64'h0166bdef9f90c4ff;
assign testcases[608] = 64'h174f0f1460b2f6f9;
assign testcases[609] = 64'h56003b83e1ffbd90;
assign testcases[610] = 64'h0e4e8fcfffecc6b0;
assign testcases[611] = 64'h087aebde7f66a0f5;
assign testcases[612] = 64'h0f08000367c8f7b2;
assign testcases[613] = 64'h07488bceffeab4a0;
assign testcases[614] = 64'h0c000b4d9ddfffd9;
assign testcases[615] = 64'h001c9fb8f5ef96d3;
assign testcases[616] = 64'hf6df76000f6fc6fd;
assign testcases[617] = 64'hfff6b033098a91f1;
assign testcases[618] = 64'h20083f8f9adff8e1;
assign testcases[619] = 64'h0f18200267baf8c3;
assign testcases[620] = 64'h220a3f8b96cdf6d0;
assign testcases[621] = 64'h0f08105085caf8e2;
assign testcases[622] = 64'h6f686005289afaf3;
assign testcases[623] = 64'he0f9df89410265c3;
assign testcases[624] = 64'h0f5fbfaf7a70c0f3;
assign testcases[625] = 64'h00174caeffabeaff;
assign testcases[626] = 64'h62100967d8ffaf69;
assign testcases[627] = 64'h61e1f9cf4f0942b0;
assign testcases[628] = 64'h00194f8ca7ecf6d3;
assign testcases[629] = 64'hfff8b250022986d6;
assign testcases[630] = 64'hef97220f6ac0f9ac;
assign testcases[631] = 64'h0d4c7dbeeffdd5a0;
assign testcases[632] = 64'h5c2b0f6fcffcf6f0;
assign testcases[633] = 64'h32a4faef6f1a0270;
assign testcases[634] = 64'h20082f6aa6fcf5b0;
assign testcases[635] = 64'hfff6a223077960c2;
assign testcases[636] = 64'h000a4f8c98defbd2;
assign testcases[637] = 64'h4f48091b7cdbf4e0;
assign testcases[638] = 64'h002b7e93c0f8fff4;
assign testcases[639] = 64'h024a2f0740b0f6fd;
assign testcases[640] = 64'h003b8fcea2e1fdcf;
assign testcases[641] = 64'h50c0f8cf4f0963e3;
assign testcases[642] = 64'h00185d88b4fafff9;
assign testcases[643] = 64'h20082f6fa9dffbf4;
assign testcases[644] = 64'h30074baaf9f3d8ef;
assign testcases[645] = 64'h00264c8f9addfde9;
assign testcases[646] = 64'h00165985c8eefffb;
assign testcases[647] = 64'h6e55083b8edffaf0;
assign testcases[648] = 64'h00062c6daeeffad9;
assign testcases[649] = 64'h0f2700277ddff9b6;
assign testcases[650] = 64'h110b7ffbf0a6fcf1;
assign testcases[651] = 64'h0a4b8ddfffdba570;
assign testcases[652] = 64'h0558acdfa8c0f7f9;
assign testcases[653] = 64'h203808115396daff;
assign testcases[654] = 64'h5f5a36097afbf6d0;
assign testcases[655] = 64'h08599ceffed79180;
assign testcases[656] = 64'h00082f7f97cdfdf9;
assign testcases[657] = 64'h645f0c6ccffcf0c3;
assign testcases[658] = 64'h00469bdf8f92e1f8;
assign testcases[659] = 64'h2039091161b5faff;
assign testcases[660] = 64'h304a1e044092d8ff;
assign testcases[661] = 64'h0174d8cfae90c0f6;
assign testcases[662] = 64'h30583f0a2274c9ff;
assign testcases[663] = 64'h0f1a246297daf5f0;
assign testcases[664] = 64'h0f3700276edffaa6;
assign testcases[665] = 64'h06488bcefff9f2d0;
assign testcases[666] = 64'h0a345382b0e0f4df;
assign testcases[667] = 64'h30084f8a92f5fef6;
assign testcases[668] = 64'h10072d6fabcefcf8;
assign testcases[669] = 64'h00184e7fbeeef9e4;
assign testcases[670] = 64'h61895f0c0360c3fa;
assign testcases[671] = 64'h0d498accffffc6b0;
assign testcases[672] = 64'h00225678aacdffff;
assign testcases[673] = 64'h100b9fa9fcbf95fa;
assign testcases[674] = 64'h0f0700388efdf587;
assign testcases[675] = 64'h1f1800278adcfeca;
assign testcases[676] = 64'ha0f4ec8f1d0560d3;
assign testcases[677] = 64'h10093f9fead7f1f8;
assign testcases[678] = 64'h40a1f6cd6f0b0371;
assign testcases[679] = 64'hb0fb98050f68d2fd;
assign testcases[680] = 64'h20482f092173c8fe;
assign testcases[681] = 64'hef99330c67c0f8be;
assign testcases[682] = 64'h340a3f7bbefdf6c0;
assign testcases[683] = 64'h0f3a333075c8f5e2;
assign testcases[684] = 64'hfff6b022088c82f0;
assign testcases[685] = 64'h0300287acdffd992;
assign testcases[686] = 64'h3f395200369bfae4;
assign testcases[687] = 64'h1f1810065adcfcc6;
assign testcases[688] = 64'h0d5dbebd83d0f9cf;
assign testcases[689] = 64'h055cacd0f4efb6f4;
assign testcases[690] = 64'hb1f5dc7f1e0650b0;
assign testcases[691] = 64'h10060c4f8bbffffb;
assign testcases[692] = 64'hd0ffaf470c6fb4c7;
assign testcases[693] = 64'habc4f6feaf5d2700;
assign testcases[694] = 64'h001a6fb8f6fffff6;
assign testcases[695] = 64'h094b8ccefff9f1d0;
assign testcases[696] = 64'hfeaf4f090160b4fb;
assign testcases[697] = 64'h0f0800458acdfbe4;
assign testcases[698] = 64'h0f4d8ecfffdba680;
assign testcases[699] = 64'h416a2d0540a3e9ff;
assign testcases[700] = 64'h90893e086ddffaa9;
assign testcases[701] = 64'h20093f8b88ccf6d4;
assign testcases[702] = 64'hef99500047a4f0fa;
assign testcases[703] = 64'h032b6f88b6ecf5d0;
assign testcases[704] = 64'h60d1f9df5f0a1384;
assign testcases[705] = 64'hffa8500149a5f8ef;
assign testcases[706] = 64'h00194f7c9adffad3;
assign testcases[707] = 64'hc0f5ec8f2c0540b3;
assign testcases[708] = 64'h5b4006388ccffbf0;
assign testcases[709] = 64'h002a6fa9b1f7fef5;
assign testcases[710] = 64'hfff7c061044894f3;
assign testcases[711] = 64'h0f3940468deff8d5;
assign testcases[712] = 64'h1f071065aafcf4b1;
assign testcases[713] = 64'h8f84500258adfff7;
assign testcases[714] = 64'he7ff98240e58b0b8;
assign testcases[715] = 64'h095cbf9b90f1fdcc;
assign testcases[716] = 64'h20051a4e9edffeea;
assign testcases[717] = 64'h71d8ff8e18009288;
assign testcases[718] = 64'h00285f8cb9fff8e1;
assign testcases[719] = 64'h06488accffdba270;
assign testcases[720] = 64'hfff7b140075bc7fb;
assign testcases[721] = 64'h2f1800367bcefad5;
assign testcases[722] = 64'h721e0094fbafb1f8;
assign testcases[723] = 64'h504c1f044083c8ff;
assign testcases[724] = 64'h737a2b0340a3e9ff;
assign testcases[725] = 64'h0f5e7e4950a0f2f1;
assign testcases[726] = 64'h705b1e0452a5e9ff;
assign testcases[727] = 64'h0f0800256bcdf8c5;
assign testcases[728] = 64'hf0faaf4f093191f5;
assign testcases[729] = 64'h10094f79bcfff9b3;
assign testcases[730] = 64'h880f107afd9fc0ff;
assign testcases[731] = 64'h05001a7bcdffc870;
assign testcases[732] = 64'h6d6118096dcff7e0;
assign testcases[733] = 64'h174f0f044081d4fb;
assign testcases[734] = 64'h0f0a022066bbfae3;
assign testcases[735] = 64'h0f4e3b4483c3f2d0;
assign testcases[736] = 64'hfff8f180013691f2;
assign testcases[737] = 64'h0f08115499fbf5d0;
assign testcases[738] = 64'hf7b651085fbad0fa;
assign testcases[739] = 64'h044689ddffca8450;
assign testcases[740] = 64'hfff5c052076bc6f4;
assign testcases[741] = 64'h30095f98c5fdfef5;
assign testcases[742] = 64'hfff7c030056ab3f3;
assign testcases[743] = 64'h7953074a9deff8f0;
assign testcases[744] = 64'h0f000348a9fcfbc5;
assign testcases[745] = 64'h1f08000548bafcb9;
assign testcases[746] = 64'h00164b8bbdfffbe5;
assign testcases[747] = 64'h120c4f8cc7d9c0f5;
assign testcases[748] = 64'h0f0a153074c7f5e0;
assign testcases[749] = 64'h10083f7f97ccfaf4;
assign testcases[750] = 64'h6b510055aaffffe5;
assign testcases[751] = 64'hef97300869c1f7b8;
assign testcases[752] = 64'hf6fd9f4d063090e3;
assign testcases[753] = 64'hc7ffcb750046b8fc;
assign testcases[754] = 64'h013467aadcffe8c0;
assign testcases[755] = 64'h001b7fa8c4fdfff4;
assign testcases[756] = 64'hfff590100a7ca2f2;
assign testcases[757] = 64'h1f0800287ccffcca;
assign testcases[758] = 64'h464f0e2470c1f8ff;
assign testcases[759] = 64'h0f2820246bcef9b5;
assign testcases[760] = 64'hc0fc97200a67d3ff;
assign testcases[761] = 64'h30070e5f89ccfef7;
assign testcases[762] = 64'h10380d064395d9ff;
assign testcases[763] = 64'h0f18004489ebf5c0;
assign testcases[764] = 64'he0ff9c310f7bd1f8;
assign testcases[765] = 64'h130f5fbef9e0a5ee;
assign testcases[766] = 64'h0d4cbc5f6760c3f1;
assign testcases[767] = 64'h0e3c7ecffffdc7a0;
assign testcases[768] = 64'h8f73260a6cdefbf0;
assign testcases[769] = 64'h0f09034388dbf5e0;
assign testcases[770] = 64'hb1f7ef8f2a0170c5;
assign testcases[771] = 64'hf7de7f1c0540b2f7;
assign testcases[772] = 64'h415a19015094e9ff;
assign testcases[773] = 64'hffb4400b78d0f8cf;
assign testcases[774] = 64'h042c8fbca3e0f8df;
assign testcases[775] = 64'h04479addffcc8660;
assign testcases[776] = 64'h00061d5e99d5f9ff;
assign testcases[777] = 64'hfff7d161014894f0;
assign testcases[778] = 64'hcf75040f7ac0f8cc;
assign testcases[779] = 64'h5f0d262057baf7c4;
assign testcases[780] = 64'hc0f9ef8c180f7dc6;
assign testcases[781] = 64'h1f073e8eefffc980;
assign testcases[782] = 64'h41094e95f8ef7a40;
assign testcases[783] = 64'h0f002e9cfadac9ed;
assign testcases[784] = 64'hc3fa9f2d0470f4f6;
assign testcases[785] = 64'h30684f0a3485d9ff;
assign testcases[786] = 64'h0c4d9f5960a4eaf8;
assign testcases[787] = 64'h20082f7f98cbf9e2;
assign testcases[788] = 64'h00185c8781e3faff;
assign testcases[789] = 64'h6f6954086acbf7f0;
assign testcases[790] = 64'h41784f093082c7fc;
assign testcases[791] = 64'h6f5604076bcefae0;
assign testcases[792] = 64'h04367aadefffd7b0;
assign testcases[793] = 64'h044488bcfffcd6a0;
assign testcases[794] = 64'h00072d6e9acfffec;
assign testcases[795] = 64'h716d1f097ddff5f0;
assign testcases[796] = 64'h20082f6f98cffed9;
assign testcases[797] = 64'h20093f8d98eef6c1;
assign testcases[798] = 64'h0f2c326098dffbf3;
assign testcases[799] = 64'h100a3f8de9c5f6fa;
assign testcases[800] = 64'h11664f0920a2f8ff;
assign testcases[801] = 64'hffe490220b6e96d0;
assign testcases[802] = 64'h000b5d94f8ff8a14;
assign testcases[803] = 64'hf4ffa950033f9ae4;
assign testcases[804] = 64'he3fbaf4f0830a1f6;
assign testcases[805] = 64'h10084d8871d2f8ff;
assign testcases[806] = 64'h0b4c9edfffca8550;
assign testcases[807] = 64'hffe772000888b1f9;
assign testcases[808] = 64'hf1feaa50030f7ed7;
assign testcases[809] = 64'h0f1800288efff8a8;
assign testcases[810] = 64'h20583f083192f7fb;
assign testcases[811] = 64'h2f18001466c6f8b6;
assign testcases[812] = 64'h0f0a152055a9faf7;
assign testcases[813] = 64'hee7f2c0450b1f7ed;
assign testcases[814] = 64'h0f08002478caf6c2;
assign testcases[815] = 64'h10073f8cbcfff8d8;
assign testcases[816] = 64'h000a4f9ba9fef7e7;
assign testcases[817] = 64'h2f130053d0b2b1f2;
assign testcases[818] = 64'h0d4e8ebefeffc890;
assign testcases[819] = 64'h0f0600468ccffbc9;
assign testcases[820] = 64'h0669cc7f6970c1f7;
assign testcases[821] = 64'h0578ed9f6a90f3f1;
assign testcases[822] = 64'hf5fcaf3e0730b0f4;
assign testcases[823] = 64'h2f49220358c9f4a0;
assign testcases[824] = 64'h0a4b8dcfffebb5a0;
assign testcases[825] = 64'hd0facc77180f6cb8;
assign testcases[826] = 64'h10464f083295eaff;
assign testcases[827] = 64'hfff7d030078a81f3;
assign testcases[828] = 64'h428f0b6470f8bdb6;
assign testcases[829] = 64'h10072f7fa9eef6c2;
assign testcases[830] = 64'h0f4e8e6c4180c3f5;
assign testcases[831] = 64'h000a5fa9e4fefff8;
assign testcases[832] = 64'h1f15055aabfcd790;
assign testcases[833] = 64'hfff7b340055ab4f5;
assign testcases[834] = 64'h6f5622046acfe8f0;
assign testcases[835] = 64'h00197fdfdca4f6ed;
assign testcases[836] = 64'h00285e8cccfff8e0;
assign testcases[837] = 64'h00375f2b4384d8fd;
assign testcases[838] = 64'h0f08102698fbf8c2;
assign testcases[839] = 64'hfff390010b8f83f1;
assign testcases[840] = 64'h22490b0350b3f9ff;
assign testcases[841] = 64'h123a0b025093d8ff;
assign testcases[842] = 64'hf3facf5f0b137092;
assign testcases[843] = 64'hfff7a213098990f5;
assign testcases[844] = 64'h807a3f093282d6fc;
assign testcases[845] = 64'h0f3902167bedf6c0;
assign testcases[846] = 64'h094b7f494092d6fa;
assign testcases[847] = 64'h0a4d9f9f6880c2f5;
assign testcases[848] = 64'h0b4e8f6f6670c2f6;
assign testcases[849] = 64'h050b1f2787f8f7c0;
assign testcases[850] = 64'hf6cf64082e94f0ff;
assign testcases[851] = 64'h3f48072a9cfff8f0;
assign testcases[852] = 64'h8f7745097bddf8f0;
assign testcases[853] = 64'h0c5dae6f6a70b8f6;
assign testcases[854] = 64'hc4fbbf4f0830a0e5;
assign testcases[855] = 64'h0f060047d8c793f8;
assign testcases[856] = 64'h0e3d7fafeffcd9b0;
assign testcases[857] = 64'hd5fc9f3e0640a0f3;
assign testcases[858] = 64'h023769abdffef7f0;
assign testcases[859] = 64'h1f09004598f9f3b0;
assign testcases[860] = 64'h0f1a142065a9f9e5;
assign testcases[861] = 64'h00083f8faad3f9dd;
assign testcases[862] = 64'h0f0800186dbffed8;
assign testcases[863] = 64'h0f18202168ccf8b4;
assign testcases[864] = 64'h90f7ff8f290082da;
assign testcases[865] = 64'h061c4f6ba9daf6f0;
assign testcases[866] = 64'h6f460b3d8edffaf0;
assign testcases[867] = 64'h0f08002066caf4d7;
assign testcases[868] = 64'hbc85300657b4f8ef;
assign testcases[869] = 64'h10098ecef9dfa8fb;
assign testcases[870] = 64'h0769bc7f6970c2f5;
assign testcases[871] = 64'h436a3f083080d4fa;
assign testcases[872] = 64'h100b5fdfcaffcffa;
assign testcases[873] = 64'h0f030047a9fafab5;
assign testcases[874] = 64'h06478acdffcc9770;
assign testcases[875] = 64'h420c7f99f6dfa4f0;
assign testcases[876] = 64'hffa740084f94f2fe;
assign testcases[877] = 64'hfff7b041045790e0;
assign testcases[878] = 64'h05498ccfffd9a280;
assign testcases[879] = 64'h0c6ebfaf5a60c2f4;
assign testcases[880] = 64'hcaaf4f0a0360d2f8;
assign testcases[881] = 64'h0f1800368cdff9b7;
assign testcases[882] = 64'h0b4b8ccefffed6a0;
assign testcases[883] = 64'h00378bcedfc6f9ff;
assign testcases[884] = 64'h00294f8dcdfdf4d0;
assign testcases[885] = 64'h00082f6dacdffbe4;
assign testcases[886] = 64'h0f39311267b9f5c0;
assign testcases[887] = 64'h10051b6b9ddfffdc;
assign testcases[888] = 64'h074a9d8f6980c3f6;
assign testcases[889] = 64'h8f77360a7ceef7e0;
assign testcases[890] = 64'h0f08201056aafbf4;
assign testcases[891] = 64'h054c9efcf4b0868f;
assign testcases[892] = 64'h10084e77abfff8d1;
assign testcases[893] = 64'h0a7ceebf7c70d8fe;
assign testcases[894] = 64'hd0f7de6f0b1481f3;
assign testcases[895] = 64'h80f4fc9f2d0561d4;
assign testcases[896] = 64'h8f6835088bfef6e0;
assign testcases[897] = 64'h00093f7e87cdfce5;
assign testcases[898] = 64'h0f043279aefff7d0;
assign testcases[899] = 64'h0f1a240054c7f4b2;
assign testcases[900] = 64'h422e0075f7cf91eb;
assign testcases[901] = 64'h20073d9bd8fefffa;
assign testcases[902] = 64'hffac50064fa7f5ef;
assign testcases[903] = 64'h07498bcdfffed7a0;
assign testcases[904] = 64'h098aec6f2e33a0f6;
assign testcases[905] = 64'hf6fd9f2c0470e3e9;
assign testcases[906] = 64'h00374f2e2561b2f3;
assign testcases[907] = 64'h0b7bec8f4d40a3f6;
assign testcases[908] = 64'h0f2830245bbffcc9;
assign testcases[909] = 64'h1f090256aaf9f2c0;
assign testcases[910] = 64'h6f67340879dcf9f0;
assign testcases[911] = 64'h0e4e9f6c5280d3f5;
assign testcases[912] = 64'hdff9d2600339a6f5;
assign testcases[913] = 64'h10062d6fabcafff8;
assign testcases[914] = 64'h6f5407297dcffaf0;
assign testcases[915] = 64'h6f5808298cfcf4b0;
assign testcases[916] = 64'h0f18102066b9f7d1;
assign testcases[917] = 64'hffa750044ba6f4fc;
assign testcases[918] = 64'h024488ccffeba480;
assign testcases[919] = 64'h0f08101569ccf9b5;
assign testcases[920] = 64'h0f1a445066b9fac6;
assign testcases[921] = 64'h095bbdffcda0e0fd;
assign testcases[922] = 64'h2f0b053487e9f4e0;
assign testcases[923] = 64'h085b9f5e3760c1f6;
assign testcases[924] = 64'h0f09123076bcfae5;
assign testcases[925] = 64'h7f66240669caf6c0;
assign testcases[926] = 64'hfff7e1400598c0f2;
assign testcases[927] = 64'h00377dbffff6c7cf;
assign testcases[928] = 64'h10061c5f8abdfce7;
assign testcases[929] = 64'h010d6fce88c0f9cf;
assign testcases[930] = 64'h0d043076bcfffac7;
assign testcases[931] = 64'hfdbf6f2d053081c5;
assign testcases[932] = 64'hf5fe9f3c0450b5fb;
assign testcases[933] = 64'hfff7b2400248a3d7;
assign testcases[934] = 64'hc0fbf266ac0f0485;
assign testcases[935] = 64'h0b5bad6f5870c2f4;
assign testcases[936] = 64'h0f1a244296e8f4c0;
assign testcases[937] = 64'hfff492200a6ea7f5;
assign testcases[938] = 64'h0459beaf5b70c3f5;
assign testcases[939] = 64'h031b4f78aeeff8f0;
assign testcases[940] = 64'ha1f6fd8f2c0460d1;
assign testcases[941] = 64'h847f0674a0fa96e5;
assign testcases[942] = 64'hf3ef77000d74e0fb;
assign testcases[943] = 64'h05488bcfffd99280;
assign testcases[944] = 64'h0f18102359bcf9d4;
assign testcases[945] = 64'h094c8edffed8a2a0;
assign testcases[946] = 64'h0f18205085c9f9f2;
assign testcases[947] = 64'hf3ffb960023895e6;
assign testcases[948] = 64'hfff6c042085ebaf9;
assign testcases[949] = 64'h1f08011066caf5c4;
assign testcases[950] = 64'hfff6b0310479a1e4;
assign testcases[951] = 64'h7f57092b9dfff8f0;
assign testcases[952] = 64'h3f58170a8bfbf4f0;
assign testcases[953] = 64'hf4fcaf4c0540a3ea;
assign testcases[954] = 64'h100a3f67acfff5e2;
assign testcases[955] = 64'h03489cc8c0f6ffbb;
assign testcases[956] = 64'h10082f7fbbfdf5c1;
assign testcases[957] = 64'h03469acf98a0e2f5;
assign testcases[958] = 64'h0b5cbeffbbb0f4ef;
assign testcases[959] = 64'h5f5520056acff9b2;
assign testcases[960] = 64'h0e5f8f4b4280d3f1;
assign testcases[961] = 64'hfff582024a84a0b0;
assign testcases[962] = 64'h3049081050a3e9ff;
assign testcases[963] = 64'h0c4c8ecffffdd7d0;
assign testcases[964] = 64'h8f67130489fcf5f0;
assign testcases[965] = 64'h085b9ebf7a80d1f3;
assign testcases[966] = 64'h42b3fabf3d0650d2;
assign testcases[967] = 64'h000a5fbeeac4f0f9;
assign testcases[968] = 64'hf8cf67022d83f0eb;
assign testcases[969] = 64'h00184f8bcffff6c4;
assign testcases[970] = 64'hef86200d69c0fabc;
assign testcases[971] = 64'hfff7b303089690f4;
assign testcases[972] = 64'h0b7bec9f6b70d6fe;
assign testcases[973] = 64'h6f4103086abdfff0;
assign testcases[974] = 64'h00185b74c6feffd9;
assign testcases[975] = 64'h0c8bfbdf7e71e0f5;
assign testcases[976] = 64'hc1f8cf5f091080d5;
assign testcases[977] = 64'h0f09122065b9f7e1;
assign testcases[978] = 64'hf4ed88170f6bc1f0;
assign testcases[979] = 64'h6048062072b6fbff;
assign testcases[980] = 64'h0a6bcdffdca88460;
assign testcases[981] = 64'h10073f7f88cdfad7;
assign testcases[982] = 64'h817c2e0540a2f8ff;
assign testcases[983] = 64'h002d8fd7f4cf96e4;
assign testcases[984] = 64'h0d4e6f5a5380d3f7;
assign testcases[985] = 64'h00061c6db9faffee;
assign testcases[986] = 64'hc0f8df7a300549a4;
assign testcases[987] = 64'hee8f3b0350b4f9ff;
assign testcases[988] = 64'hfff58100097aa0e4;
assign testcases[989] = 64'h744c0a2270c2f9ff;
assign testcases[990] = 64'hf7ffc7700043a3b5;
assign testcases[991] = 64'h0c4c8ddfffc68055;
assign testcases[992] = 64'h0f3940357bcef9d6;
assign testcases[993] = 64'h5248071060a4eaff;
assign testcases[994] = 64'h20574f0b0264b7fc;
assign testcases[995] = 64'h2f15001a87f5b3f3;
assign testcases[996] = 64'h00071d5f8bcafae4;
assign testcases[997] = 64'hfff5c140056ab2f1;
assign testcases[998] = 64'hff99400b5ea2f1d9;
assign testcases[999] = 64'h0f2700378dfff9d8;



pendigits_tnn1_tnnpar dut (.features(features),.prediction(prediction));

integer i,j;
initial begin
    features = testcases[0];
    for(i=0;i<TEST_CNT;i=i+1) begin
        features = testcases[i];
        #period
        $display("%h",features);
        $display("%b",dut.hidden);
        for(j=0;j<CLASS_CNT;j=j+1) begin
            $write("%d ,",dut.scores[j]);
        end
        $display("");
        $display("%d",prediction);
    end
end

endmodule
