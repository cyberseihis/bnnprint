













module pendigits_bnn1_bnnroperm #(

parameter FEAT_CNT = 16,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 10,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 640'b1110000011011010010100011111000011001010000111010100111000011011111010010101101001101010010100111001001000111101010010100001101100010110101111011010010000110111000101101110110110110001000001110100001111101100010111111100000110111010111001010101101001100011000000000010111101010001111100001011000000101011111110111101000001001011111110001110111110000101011010111111100001001010011000101011011011011001010100000101100110110101000010011011110100100011010010111010010000000111000010111011001011110101010011010001101010100101110010001001010101011000101001010001111000000101001110001010111110110001000000110101001011011010111101010010101101000010 ;
  localparam Weights1 = 400'b0011000010000110000111010101111000001010100010101101101000110110101110101100001011111001000010000101100111000011101010100011010011110000101000001011010010001000101101000100001010101110100111100011101000011001001011010001010000111101000000110101111011100100010110111100011111111100111111101010100101001001110000010000010011101010101011011101111101001010000001100000111000010110000101001011010011101101 ;

  romesh_seq #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
