
















module Har_bnn1_bnnpaar #(

parameter FEAT_CNT = 12,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 4448'h0064008700560086004f00790068007800520077005900760049007500490074004a007200630071005c00700044006f0045006e0061006d0042006c0045006b003c006a0055006900570067005a0066003b00650046006200420060004e005f003c005e0054005d0046005b003b00580036005400220053001d0053003f0052003e0051002b0051004b0050002b00500047004f004d004e0040004d004a004c0043004c001e004b003b00480024004800330047002a004400340043003c00420032004100330040002e00400031003d001c003a00340039002e003800210038002900370027003700280036002c003500260035001d0035002900300026002f0027002d0020002d0023002c0019002b0028002a0024002a001b00280023002500200025001c002500210022001b002200180020001e001f001f0041002a003f001a003e0018003d0032003a0030003900360038002e003700280035001d00310024002f002d002e0021002d0029002b001a002b0026002a002500280020002400310034002200330018003200270030001d002f00230029001c0027001b00250019002400180019001c002c001b002600030015001e0023001a002200110014001c001e00040016000e0012000a0010000500080002000600000001001d0020001a001b0009000f0007000b00180021001300170001000c000c000d0019001f00070017000800110004000a0006000e00030009000b00130002001200100016000f0015000500140000000d ;
localparam YMAP = 640'h00a1007c008800970081008e0095008a00930083009800850084008b009f008f0080008c007b009c009100940090009b007f0089007d0073009a009e008d007a009d007e00a2009200960099008200a0;
localparam ADDCNT = $bits(PAAR0) / 32;
localparam FULLCNT = ADDCNT + (FEAT_CNT * 2);
localparam Weights1 = 240'b111001111101100000101111100101100010100011010110111111001010010101011010011101001110011111011110001101011100001000101010010101000110011010101101110010110100110101111111011000000011000110001111110000010111001001000101000010011100001111000100 ;
localparam WIDTH = 320'h06060607070607070707070807070707070707070707070707080707070707070707070708070707;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[FEAT_CNT+i] = -feature_array[i];
endgenerate

integer j;
generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam op1 = PAAR0[i*32+:16];
    localparam op2 = PAAR0[i*32+16+:16];
    localparam nodeloc = (2 * FEAT_CNT) + i;
    assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    assign hidden[i] = node[YMAP[i*16+:16]] >= 0;
end
endgenerate

/* initial begin */
/*     #10 */
/*     for(j=0;j<FULLCNT;j=j+1) */
/*         $display("%d | %d", j, node[j]); */
/* end */

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wneur[j])
            tmpscore = tmpscore + hidden[j];
        else 
            tmpscore = tmpscore + hidden_n[j];
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = tmpscore;
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
