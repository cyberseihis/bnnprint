












module winered_bnn1_bnnshift #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 440'b11111100010011001010011010011110111010001111101010001001111001011011101001000000110011100011010111100110111100111111101101011100001111000001110100111011000001111011100110100100011001101101101000100110101111010101101100111100100010011000000001011111111000110111000111001011011000010000000001010111011110110010000011100101101110001100011001101011101101101001100011011010011000000011001111000110101100001000011100101000111100001111001001111000 ;
  localparam Weights1 = 240'b101011110101010111101111010101000101111001101110110011111110010011110100100011101000101011111101111001010101001011000101101011100011011000100010000100100000001111000110100000011011100000011101001111010010001011110000001101110000010000111001 ;

  seq_bnn #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
