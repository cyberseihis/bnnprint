











module winewhite_tnn1_tnnseq #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnn #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(440'b10000000101000101101000100000010000101100001100001001000000000010100000000010110000010000000000011100000001010000000010000000011110000001010010100010010010000111010100000001001100011011000111101100010100001101110000010010011000101000001100000000101010010001000000100101010010000110000010101001010000001010100010001010010010010010000000111000101011110010100011001111011000000011111110101011001110000000000100000100001011100100000000010001000),
  .MASK(440'b11000000101101111111010101111010100101100011100001101000001010010101100101010111100010000010000011100110101010110000010110011011111000111011011111010110111011111011110000001001110111011100111111101110101101101110000111011011001111011001110010101101010010101001101101101010110111110010110101101111011011011100011001110010010111010010110111001101011110010110011001111111111000111111111101011001110110011000100010100001011100100000001110011001),
  .NONZERO_CNT(640'h07030606090603050506090105030508080807070707060904080506080407070707040706080706),
  .SPARSE_VALS2(79'b0100000010110010011000100000110000101111111100111011000110111010101011011001010),  // Bits of not-zeroes
  .COL_INDICES(632'h2625232221201e1b1817141211100d0c0605040201211f17100d0b211c1615100c0825211f1817100f0125242119181412092625221f1e1c1817161413100b0a07261c171412100f0b0a0907060401), // Column of non-zeros
  .ROW_PTRS(64'h4f3a342d251d0e00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
