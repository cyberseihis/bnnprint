











module gasId_tnn1_tnnseq #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnn #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(5120'b10000000010010000101001110000000001100011001000000101000010100111000000000010000100000110100100000010001000000000000000010000000011000000001100110100000011100001000000101001001011110011010000110100000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000100000001000000000000001000000100010011100111000101011100000011001001110100000010010100010000110000000000100001000000001001010001010111010000100010001100000010101101000101011101000010001001100111001100011100110001010000001110101110000000000000001000000010000000000000000001001000000000000000000000001000000000000000011000000000000000000000000001000000010100000000110001000000000010010000000001110001000010011100110010010000000010001110001100101001000000000000000000011000101100110001101111000100001100010100010100100000100000000010000000101000011000000100010000000000000000000000000000010001000000000000000001000000000000001000000000000100000000000100001000000000000000000100010000000000010001000000001010000000111100010000100111001010100100000001100001110001001010010000110001001011000110101000001100001001110000100011010101010000011000001100000010100010101000001110010101000100000000000000000000001000100000000100000000000000000000000000000000000000000001000000000000000000000010000000100001100000010000000000010000000001000000000000000001000010000000000000000100100001000011001110000000110000011110001001000111101000110000000010101010101000010000000100011001000000010000000000010010000000010001000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000100000001000000010000111001000000000100110000000000000000000000000000010000100001100001001100000110000000010000111010000100000100101000101100000101000000000100000010011100000100000001000110000000010100000010010000100000000010000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000010000000110010000000000000000000010010000000100001010000000000001001010000001000000000000100000011010000000100010001010100001001001100010101010000001100000100000100100000000100000001101000100000000000010000000000000000000000000100001000000000000000000000100000000000010000000000000000000000000000000000000000000000001000000000000000000000000000010000001000000000011000000000000000000000000000000010001100000000000001000000000000000000010001000000000010010101010110000010100000000000000000001001100100010000001110000000000000000001000000000000100000110000000000010000000000000000000000000000000000110010000000000000000000000000000000001000000001101011000110011000000000110010100001000111000000001001101100010011100110000000011010000101000111000000011100001000000001101000000100011000000001110010100100000110101001010011100000000111001000000010000000000000100000000000000000000010000000010000100000000000000000000000000000100000000100000000000000000100000010110000011010000101001111000100001100001110011001100000000100010101010000110000111001000110000000010001010100000010000011100100011000000001010101010000001000001011001001101000010100011100000000110010001000000000000100000000000000000000000000000010000100000000000000100000000000000000000000000000000000000000000000001000001110001000111001000011000000000000000101111010100011001100001101000000011001010010100011010100010000110100000000000101011101101000010101000101010000000011000000010000100011100100001100000010000001000000001100000000000000000000100000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000011010000000000000000000001000110001000010001000100010000000100010000100011000000010010100000000001010001010100000100000100010000010001100001100000000001100001000010001001001110000110100000000010000000000000000000000000000000000000000000000010000000000000011000000000100000000000000000000000000000000110000000100010000000100001000000100001110000000000010100000000100010000011000010001000100001000110000000110000001111001000100011000110011000000001000101010000001010001101000100101100110101010101100010100010000000010000111000000011000000000000000000000000000000000010000000000000000000000010001100000001000000000000000000000000101000110000001000100010001000001000000000000000000000001010000000101000100010001000000000100000000100000011010011001000100001000110000100010001010100000110100001010101001011001101010101011000101000100000000000000001000000100100000000000000001000001000000000000000000000000000000000100010000000000000010000000000000000000001101000001010000000111000010100010101010100001000110001000101010000000010000001001000010000000100000100000100000100000101000010001100010001010101000000110000110011101100010001011101010110000011000000000000000000000000000000000000000000000000001000000001000100000000000000000000000001100000000000100000000000000000000000000010000000100000001010000000000000000100000010000100010010010101100001100000000000000100000000000001010001000000000001010100101001001101010101011000001000001101010001100000010100010101000000110000000000110000000000000000000000000100000010000001000000010000000000000000000000000010000000000000000000000000000001000000),
  .MASK(5120'b10000100010110001101011110101010101111011001001010111001010100111010010000011001100000110101100100010011000011000100000010110000111000000101101110100000011101001111000111011001011111011110010110100100100000000001000000100000000000100100000000000010000000000000000100000000000000000000000000100000001000100000010001000000110011011111111010101111111111011011101111100101110110101010010111010100000101001111010011101110111011111111110100111001111101011111111011101111111111010101101101111101101111100111011111011101111111110000001000001001000000010000000000000000001001000000000000001000000001100000001000100011000000000000000000000010001000001010101001100111001110000011011010110000101110001110010111111111011010000011010011110001111111001001100100000010001111000111110111111101111010100011111110101011100100101101010000011110000101101111010100110010000000000000000000000010000010001000000000000000001000100000001001000000000000100000000001100001000001000000100010100010010000000011101000000001011100001111100111100110111111011110100100011110101110001111110010011111101101011011111111000001110001101110100100011111101010010011101011110111111110110111000111110111101000100000000000000000000001000100000000100010000000000010000000000000000000000000001000000000000000000000010000000100001100011010110110001011000001101010000000000010001100010000010000000000100101001011111111111111010110101011110011011011111111011111001000111111111101011010010100100011001000000010000001000110011100000010001000000000001000000000010001000000000000000000000000010000000000100000000000000010000000000000000000000100000000000110000010100100011000010010000111101000000000100110000000000000000000100100000010111101101111101101101111110010000111100111111111111010101111111111101110111011100010100100010011100000100001001001110001000010100000010010000100000010010000000000001000000001000000000000000000100000000000000000000000100000000000100100000000100110001000110010010000010010001000010010001000100101010010000000001001010000101000000000000100000011010000001100010011110101001001111110010111110011101100000100001100100010000100100001111010100001000000011000000101000000000000100100001000000010000000001000100000000110010000000000001000000000000000000000000000000000001001000000000000000101000000010000001000000000011000110010000000000100000000000010001100000000000001000000011000000000010001100000101010110111110111011010100100101000000000111001101100010010101110000000000000000001000000000000111001110000000000110000000000000000000001100000000000110010000000000100000000000100000000001100110011111111100111011010101010111110111111011111010001001111111100111111100110000101111111001111000111101100111111001000100011111100101101011010110011111111100101001111101011010111101011101111111010110111000001000010100000000110000000000010000000010000100000000000000000000000000000100000000100000010000000000100000010110100111111011111101111101101111111011110111111101110011100111111011010110100111011011110001001010011111100011010000011101100111110110111011101010001101001011011001011111000111110011110000110111111001000100000000100000000000000000010000000100010000101000000000000100010010000000000000000000010000000000000011001001000001110011010111011011011001100000000100111111010111011001101001101110110111011011010110111110101010100110111000010101101111101101010011101101101111001111011000000010100101011110101001100100010000001000000001100000001000000000000100000000000000000000000000001100000000000100100010000100000000000110010000000000000000000000100010100100011010100010001011000100001100110001010010101110100011000000110010010100011001000010011100000010101011001010110000101000110010000111011100111100001001101110001011010101011001111100110100000000010000000000000000000000110000000000000000000000010000000000000011000001000100000000000000000100000000000000110000001100011100000100001010101110001111101000011111111001010100010110111010010011001101011011110111001110001011111111001110111101110111011100111001111010011101011011101000101111110110111010111111110101011000000010000111000000011000001000000000000100000000000000010000000000000000000000010001100000001000000000000001000000000111010111100001100101011011000101011010000001000110010101010001111101010100110011100101110101110010100111111011011001101101011011110111101110011110101111110110101010101011111101101111101111111111010110000000100100001000000100110010010001000001000001000100000100000000101000000000000100010000000000000010000000000000000000001111000011010100100111011110111111101010100001010111001100101011000011110000001001011010000000110000100000100110100000101000010011100011001110111000110111001111011111100011001011111011111011011000100000000000000000000000000000000000000000000001000000001000100000000010000000000000001100000000000100000000000000000000000000010001000100011011010110000111000000100000010000110011010111111101111100000000000110100000100100001011001001000000001110101111111101111111111111001101000111101011001110010011100010111000111111001000000110000000000000000010000100100000010000001000000010000000000000010000000000010000000000001001000000000001001000000),
  .NONZERO_CNT(640'h3427422822283d33363239252b30332a24333d3328233544252e372f1f3d392639323e2d2d261429),
  .SPARSE_VALS2(58'b1000100000101101101100001111000000101101100010010010010110),  // Bits of not-zeroes
  .COL_INDICES(464'h2419161514110d06040327241816150c0805041d110c2322201d1c1a19110c090600251f1c1513100d0b0a0908002722201f1d1a16130e0a0802), // Column of non-zeros
  .ROW_PTRS(56'h3a302724180c00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
