











module cardio_tnn1_tnndirect #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnndirect #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(760'b1000001000111100001100110000100110000010000000000100010100100000000110101010110100000000000000100001000000001000110000110100000100001000110000001010101010001011011101100100000000101101001110000001000000000000001010000000001000100000101011100100010001100010000000101000000000001000010000010000010010001011000100010000000000001000000000000000100001101001000001000000001010011010011010000000011000101000010100010000101010000000000010010101000001010000011000000000001010000000000000000001011000000001011100000000010101010000001001000100000000010110101000000000010010100100001000000001000010001010001000000000000010000100010000100010100000001001000000010000100100101000101001000100000001010100000001100000001001000000010001101101100010000000001001000100000000110110),
  .MASK(760'b1100101000111101011111110000101110101011000000110100111100100000011110111010111100110000010010100001100000101010111100111101000110111100110000101110111011111111111101111100101010101101011111111111100000001000101011000010001100110000111011110110010101100011101000101010000010101000010010010001011011001011000110010010011010101000000000101000100011101001000101011000011011111110011011100100111110111100010100010101101010000000100111110101001001011010111010100001001111110101110000000001011100000011011100110010111111011000001001001110000110010110101001010010011111100110101000100001110111011110011001100100000010010110110100110110111100001001001011010100110110111101101111110101000101110101010001110101011001010110010001111101100110000101001101100100000000110110),
  .NONZERO_CNT(640'h0b0b090909070c0a110c09080a0906090804090b0d08080a0b040d08080b0a070b090c0c0a0a0807),
  .SPARSE_VALS2(39'b101110010111100011111111011101111110001),  // Bits of not-zeroes
  .COL_INDICES(312'h26211f1b130f0d0b080705040225211e1c1b0f0c090706050201252421201c1b1a18110c0a0301), // Column of non-zeros
  .ROW_PTRS(32'h271a0d00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
