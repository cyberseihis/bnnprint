












module winequality_white_bs #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 5


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 440'b01011011001001010110011000111111100001101110011110111101111010000011000010100110111100010000110010110011100101010111010001001000111000101011010101001110010111011110101100111011111000110011011010110110011111001000001111001101001001101000010110100001111111101110001001001000111100001010010111011000101010001111011111100101110010110001011100100001001001110010100011000000000001001011010100011010101110001001110001001010111111100000111001011000 ;
  localparam Weights1 = 280'b0110101101111010110110010101001100000000111001110111011111111000110100011011000011101011011100101111000011010111101100001100101101000010001100000101011110110000111010110111001011111000110101111101100011101011011100101111110011000111101100011110001101010011010011001100000001110011 ;

  seq_bnn #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
