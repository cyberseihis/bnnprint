











module cardio_tnn1_tnnseq #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnn #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(760'b0011110101000000000000001000000001110001101000000000010001101010101110111010110011001000000010000001100000000010000000000010000000000100011001001110001010001100101001010111000000010000000000010000000010000000000000001110100000011001111010110000011000011000100000000000001000000011000000000010001000001000100000011000110100110000000100100101100001010011000010010001011101111000000101000001001100000010000010000000001100100000100100000000000000000000000100000000100100100011010000000100010000100001100001000001000100000001000000011000010000001000000001000100000010001000000001001010010000010001111000100000000000000100000001010010100010010010011000000000100000100000101000000000000001011110100001000000001000001000000110001000000101001000000100000000000100010111),
  .MASK(760'b0011111101000100000001011100111001110001111111110111110111111110101110111110111111101000000011010001100100000011110101000011011101101101111101001110001110101111101011010111010000010001000111110100110011010100010000011110111100011001111110110000011010011110111110001000001010000011010100010110001111011010101100011010111100111100011100110111100101010011000010010001011111111101110111001011101111001110000010011010011100111000111100010000110000100100001100011000100100100011010100000110110100100001110001001101010101010001010110011000010000011000000101110110000010101010110101001010110100011101111000110001111100111101000001010010111110010010011010100000100000110100101001010001001011011110100001001001001000001111010111111000000111101100000100000110010111010111),
  .NONZERO_CNT(640'h07080a0a0c0c090b070a0b08080d040b0a08080d0b0904080906090a08090c110a0c070909090b0b),
  .SPARSE_VALS2(39'b101110010111100011111111011101111110001),  // Bits of not-zeroes
  .COL_INDICES(312'h26211f1b130f0d0b080705040225211e1c1b0f0c090706050201252421201c1b1a18110c0a0301), // Column of non-zeros
  .ROW_PTRS(32'h271a0d00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
