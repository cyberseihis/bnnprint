











module winequality_red_ts #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnn #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(440'b00000000010001000100001100110110101110100000110011001011000000000000110000000010100011011100011001100001101010101000000000000000110000100000010001100001100010100001100010000000000000101001010000001010100001000000011000110101111000001001000101010100100001110110001000000100011000110000000100000010101110001000100100000011010100000000010000100001001000101000000010000100001000000100101000000000010100000000000101011100101100100101001011000000),
  .MASK(440'b11000101110001000101111100110110111110101010111011111111100000110110110110001110100011011111111011101001101111101111000111000010110000101000010111100001110110101011100110000010011001111011010001001110111111010101111011110101111000101001100111010111101101110111001101011110011100111000110100111010101110001010101110011011010111000000010110110101111000101011001110101110101011010101111010101111011100010101100111011100111101101111001111100001),
  .NONZERO_CNT(640'h09060405080804070806050606080704070707070407060808060a05050608050807060806020707),
  .SPARSE_VALS2(71'b11111010010011110001001011010000111010010110011001101111011010010001010),  // Bits of not-zeroes
  .COL_INDICES(568'h2523211e190e0d0c08060400252421201f1d1916140f0e0c0b070302010027222120170c06012321190e0d0c0908040100231d1c0d0b0a0905271e1d1c1a171612110c04030200), // Column of non-zeros
  .ROW_PTRS(56'h473b2921160e00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
