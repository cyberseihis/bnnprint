module doublesum (
input [30:0] a1,
input [30:0] a2,
input [30:0] a3,
input [30:0] a4,
input [30:0] a5,
input [30:0] a6,
input [30:0] a7,
input [30:0] a8,
input [30:0] a9,
input [30:0] a10,
input [30:0] a11,
input [30:0] a12,
input [30:0] a13,
input [30:0] a14,
input [30:0] a15,
input [30:0] a16,
input [30:0] a17,
input [30:0] a18,
input [30:0] a19,
input [30:0] a20,
input [30:0] a21,
input [30:0] a22,
input [30:0] a23,
input [30:0] a24,
input [30:0] a25,
input [30:0] b1,
input [30:0] b2,
input [30:0] b3,
input [30:0] b4,
input [30:0] b5,
input [30:0] b6,
input [30:0] b7,
input [30:0] b8,
input [30:0] b9,
input [30:0] b10,
input [30:0] b11,
input [30:0] b12,
input [30:0] b13,
input [30:0] b14,
input [30:0] b15,
input [30:0] b16,
input [30:0] b17,
input [30:0] b18,
input [30:0] b19,
input [30:0] b20,
input [30:0] b21,
input [30:0] b22,
input [30:0] b23,
input [30:0] b24,
input [30:0] b25,
output [35:0] outa,
output [35:0] outb
);

assign outa = a1+ a2+ a3+ a4+ a5+ a6+ a7+ a8+ a9+ a10+ a11+ a12+ a13+ a14+ a15+ a16+ a17+ a18+ a19+ a20+ a21+ a22+ a23+ a24+ a25;
assign outb = b1+ b2+ b3+ b4+ b5+ b6+ b7+ b8+ b9+ b10+ b11+ b12+ b13+ b14+ b15+ b16+ b17+ b18+ b19+ b20+ b21+ b22+ b23+ b24+ b25;

endmodule
