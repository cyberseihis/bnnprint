












module winered_bs #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 440'b00011110010011110000111100010100111000010000110101100011110011000000011001011011000110010110110111010110011000110001110110100111000001001101111011101010000000001000011011010011100011101100011111111010000000011001000100111100110110101011110101100100010110110110011000100101100111011110000011011100101110000011110000111010110111111100111101100111101011000111001100000010010111011010011110010001010111110001011101111001011001010011001000111111 ;
  localparam Weights1 = 240'b100111000010000011101100000011110100010010111100101110000001110110000001011000111100000001001000010001000110110001110101101000110100101010100111101111110101000101110001001011110010011111110011011101100111101000101010111101111010101011110101 ;

  seq_bnn #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
