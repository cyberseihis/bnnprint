











module Har_tnn1_tnnseq #(

parameter FEAT_CNT = 12,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnn #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(480'b000001000000000110011100000100101100000110001100000001001100100001100000000000010000100000001011000101000001011001100010010000001100000000011011000001001011001110100110000100011010000001111000001100000010001000100111001010000101000010110001000000000001000001001100000100110010001001001110001000100001000000010000000000001001000011101011000001011000110001011010000000010000010010000000010010001110100000011111100010100000000010100010100000111000000011100000000010110110001000100000),
  .MASK(480'b110011110011001110011111101110101101110110011101000001001101100111101011000100011010100101011011111101110011011011111011110010001101000101011111000001001111001110100110101101111110100001111010101100110010111010101111001010100101001010110001001100111001000001001100101101111010101011011111101011101101000000010100100011011001011111101111001011011110111111011011001000110110011010001000010011111110101000011111111011110001101010100111110000111111111011110010100011111111001010101001),
  .NONZERO_CNT(640'h08040606080809080806080605070907070604060a0606060606080705070a050b0607070702070a),
  .SPARSE_VALS2(89'b10010110011111001000011111001110110110101011011001101110001000101101101100100001101100111),  // Bits of not-zeroes
  .COL_INDICES(712'h272623201d1b1a1712110d0b03002623201f1d19120e0c0b0805042622201f1d18151211100b04010021201b1a1918161512110d0a060100242322211f1d18161412100e0c0b0a06052422201e1c1a1918161411100e0d0a06), // Column of non-zeros
  .ROW_PTRS(56'h594b3e30211000) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
