`timescale 1us/1ns





module tbcardio_tnn1_tnnseq #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000




)();
  reg [FEAT_BITS*FEAT_CNT-1:0] data;
  wire [FEAT_BITS*FEAT_CNT-1:0] testcases [TEST_CNT-1:0];
  reg rst;
  reg clk;
  parameter Nsperiod=50000;
  localparam period=Nsperiod/500;
  localparam halfT=period/2;


assign testcases[0] = 76'h4000d18100621208964;
assign testcases[1] = 76'h8203140320b3a52a991;
assign testcases[2] = 76'h8103140420b3a42a991;
assign testcases[3] = 76'h8104150720a07a0a991;
assign testcases[4] = 76'h8203150600a0780a991;
assign testcases[5] = 76'h81073d0098d0b45254a;
assign testcases[6] = 76'h81064e0068d0b55154d;
assign testcases[7] = 76'h5000f11500621008770;
assign testcases[8] = 76'h5001f11400621008770;
assign testcases[9] = 76'h5002f01300621108770;
assign testcases[10] = 76'hd001b42910b1920bbb1;
assign testcases[11] = 76'hd001b41910b1940bbb1;
assign testcases[12] = 76'h7224330420664409990;
assign testcases[13] = 76'h744333021083520a991;
assign testcases[14] = 76'h74e325026492760a895;
assign testcases[15] = 76'h7282150334927309883;
assign testcases[16] = 76'h7282340330b0840a894;
assign testcases[17] = 76'h7171150434927409883;
assign testcases[18] = 76'h7193240334915509782;
assign testcases[19] = 76'h74f4440254a28529882;
assign testcases[20] = 76'h709344032cb18c09568;
assign testcases[21] = 76'h7281340224c1a809882;
assign testcases[22] = 76'h7061550128d1ba22449;
assign testcases[23] = 76'h7000f10200191008770;
assign testcases[24] = 76'h7001f0e100191009880;
assign testcases[25] = 76'h5000f0d1001a1108770;
assign testcases[26] = 76'h5000f022002b3108870;
assign testcases[27] = 76'h5000f0c1001a1008770;
assign testcases[28] = 76'h80514a03a4c0a629784;
assign testcases[29] = 76'h80203e0280d0a909665;
assign testcases[30] = 76'h80413a04c0d0b809773;
assign testcases[31] = 76'h80222f02a0d0b908664;
assign testcases[32] = 76'h8021460570d0aa29782;
assign testcases[33] = 76'h4631380710b18c08771;
assign testcases[34] = 76'h4421370410b08829871;
assign testcases[35] = 76'h4334380800d0aa08771;
assign testcases[36] = 76'h3434280630b08807661;
assign testcases[37] = 76'h2202370520c09707661;
assign testcases[38] = 76'h3312280610c09707661;
assign testcases[39] = 76'h3623350400b08607761;
assign testcases[40] = 76'h2626350410914627761;
assign testcases[41] = 76'h2214350400b18507761;
assign testcases[42] = 76'h3112630400814508771;
assign testcases[43] = 76'h3203640400d0ac28771;
assign testcases[44] = 76'h50012a0540d0b607661;
assign testcases[45] = 76'h50012b0540d0b707661;
assign testcases[46] = 76'h50031b0720d0ac08771;
assign testcases[47] = 76'h51032b0720d0aa08772;
assign testcases[48] = 76'h51032f0540d0b609774;
assign testcases[49] = 76'hf406340510b4a60eee1;
assign testcases[50] = 76'hf2044304005ea40eee1;
assign testcases[51] = 76'hf006790750d0b62bab4;
assign testcases[52] = 76'hf0065c0164d0b707996;
assign testcases[53] = 76'hd000a172103c520ccb0;
assign testcases[54] = 76'hc000c0c2001d430bbb0;
assign testcases[55] = 76'hd000a29420b19b2bbb0;
assign testcases[56] = 76'hd000a39410b19b2bbb0;
assign testcases[57] = 76'hc0036172001e610ccc0;
assign testcases[58] = 76'hc0036152002e610ccb0;
assign testcases[59] = 76'hb30342020094840bcb0;
assign testcases[60] = 76'hc2036232004c840ccb0;
assign testcases[61] = 76'hc2026142002e720ccb0;
assign testcases[62] = 76'hb0013304002c500bba0;
assign testcases[63] = 76'h9103330400a49a0aa90;
assign testcases[64] = 76'ha10333040094890aaa0;
assign testcases[65] = 76'hd0026172001e510ccb0;
assign testcases[66] = 76'h910272440095883dcc0;
assign testcases[67] = 76'ha3025203005a820ccb0;
assign testcases[68] = 76'ha3025203005a820ccb0;
assign testcases[69] = 76'hb0047104003c640dcc0;
assign testcases[70] = 76'hb1037104002d630dcc0;
assign testcases[71] = 76'ha60293050093700bba1;
assign testcases[72] = 76'ha40093040093720bba1;
assign testcases[73] = 76'ha50394060093720bba1;
assign testcases[74] = 76'ha70593050093730cbb1;
assign testcases[75] = 76'he001b2040084620ccc0;
assign testcases[76] = 76'hd001a213002d600ccb0;
assign testcases[77] = 76'hc201530400a1732bbb1;
assign testcases[78] = 76'hc101540700a1752bbb1;
assign testcases[79] = 76'hc202540700c1a40bbb1;
assign testcases[80] = 76'hc001540800a1642bbb1;
assign testcases[81] = 76'hc101630600c1a82bbb0;
assign testcases[82] = 76'hc001620500c1a72bbb0;
assign testcases[83] = 76'hc401730000a2740ccc1;
assign testcases[84] = 76'hc611620400b2940ddd1;
assign testcases[85] = 76'hc711620000a3940ddd1;
assign testcases[86] = 76'hc301640700a0640cbb1;
assign testcases[87] = 76'ha010630410c09409990;
assign testcases[88] = 76'ha000b15400a3940bba0;
assign testcases[89] = 76'ha100850220d0bb6b9a3;
assign testcases[90] = 76'ha101b052002c610dcc1;
assign testcases[91] = 76'hc000c0c2001d440bbb0;
assign testcases[92] = 76'hc000c0c2001d420bbb0;
assign testcases[93] = 76'hc000c0d1002b430bbb0;
assign testcases[94] = 76'hc001d0d1001d400bbb0;
assign testcases[95] = 76'hc000a113002c510bbb0;
assign testcases[96] = 76'hc000b053003a532bbb0;
assign testcases[97] = 76'hc000a1921074530ccb0;
assign testcases[98] = 76'hc000a172103c520ccb0;
assign testcases[99] = 76'h640114020087a729980;
assign testcases[100] = 76'h6201341420836309881;
assign testcases[101] = 76'h6401330510574539880;
assign testcases[102] = 76'h6301330500734409980;
assign testcases[103] = 76'h61004203002a3009880;
assign testcases[104] = 76'h6100240500734429880;
assign testcases[105] = 76'h6312260550b19428771;
assign testcases[106] = 76'h6010290440d0a628661;
assign testcases[107] = 76'h6202240410938708871;
assign testcases[108] = 76'h6313250240c2a728871;
assign testcases[109] = 76'h6000330600543428870;
assign testcases[110] = 76'h6211250140b4b909871;
assign testcases[111] = 76'h7401540400a4a90a990;
assign testcases[112] = 76'h720253030087a50a990;
assign testcases[113] = 76'h7001620400596429980;
assign testcases[114] = 76'h73042c0080d0ac2a785;
assign testcases[115] = 76'h70022b0070c09639664;
assign testcases[116] = 76'h50023a0614d0a728557;
assign testcases[117] = 76'h5203420250574308770;
assign testcases[118] = 76'h5102420140564308770;
assign testcases[119] = 76'h5102330130564308770;
assign testcases[120] = 76'h5004725250b19c39771;
assign testcases[121] = 76'h5002816130846608770;
assign testcases[122] = 76'h5002723140713728771;
assign testcases[123] = 76'h5202430120c2b829772;
assign testcases[124] = 76'h5003330134722327661;
assign testcases[125] = 76'hf003b0330085700ddd0;
assign testcases[126] = 76'hf002c042001f600ddd0;
assign testcases[127] = 76'hf001b1140085700ddd0;
assign testcases[128] = 76'hf001b022001f600ddd0;
assign testcases[129] = 76'hf00091630084730ddd0;
assign testcases[130] = 76'hf0009172001f700ddd0;
assign testcases[131] = 76'hf00091530084610ddd0;
assign testcases[132] = 76'hf000a1a1001f700ded0;
assign testcases[133] = 76'hf107a013004c840ddd0;
assign testcases[134] = 76'hf104a102004c840ddd0;
assign testcases[135] = 76'hf004c023002f700ddd0;
assign testcases[136] = 76'hf104a102004c840ddd0;
assign testcases[137] = 76'hf003c032002e700ddd0;
assign testcases[138] = 76'hf106a113003e900dee0;
assign testcases[139] = 76'hf104a123004e920dfe0;
assign testcases[140] = 76'hf001a103002f810eed0;
assign testcases[141] = 76'he201740810d0a9fccc2;
assign testcases[142] = 76'he00182040086840ddd0;
assign testcases[143] = 76'he101740b00d0a78ccc1;
assign testcases[144] = 76'hb402821500b1890bba1;
assign testcases[145] = 76'hb30182010093840bbb0;
assign testcases[146] = 76'hb10182260093772bba0;
assign testcases[147] = 76'hd10282160093740bcb0;
assign testcases[148] = 76'hd10082230084742ccb0;
assign testcases[149] = 76'hc1039133004a662ccb0;
assign testcases[150] = 76'hc001a143004a640ccb0;
assign testcases[151] = 76'hc0019123004a540bcb0;
assign testcases[152] = 76'ha403640310b07b2cbb2;
assign testcases[153] = 76'h620343040079b308981;
assign testcases[154] = 76'h600252050079b408870;
assign testcases[155] = 76'h5103622300394208870;
assign testcases[156] = 76'h5103612300293208870;
assign testcases[157] = 76'h51036223002a3108870;
assign testcases[158] = 76'h55055221003a3108870;
assign testcases[159] = 76'h53034211003a4208870;
assign testcases[160] = 76'h52035231003a4108870;
assign testcases[161] = 76'h52035221003a4108870;
assign testcases[162] = 76'h5204422310724208770;
assign testcases[163] = 76'h5203422300654228870;
assign testcases[164] = 76'h5202422300553408870;
assign testcases[165] = 76'h8201970d10b1910a991;
assign testcases[166] = 76'h8101980f00b1910a991;
assign testcases[167] = 76'h8101c31800c1a20a990;
assign testcases[168] = 76'h8101c20500b3a50a990;
assign testcases[169] = 76'h3101717200462408770;
assign testcases[170] = 76'h3002714210611508760;
assign testcases[171] = 76'h3001815200191108770;
assign testcases[172] = 76'h4102430310846328770;
assign testcases[173] = 76'h4101430400846338770;
assign testcases[174] = 76'h4101431400846508770;
assign testcases[175] = 76'h4202430300c1a608870;
assign testcases[176] = 76'h4001520400814408870;
assign testcases[177] = 76'h4503440310b3a809991;
assign testcases[178] = 76'h4102330410563308770;
assign testcases[179] = 76'h4401440200c1aa0a991;
assign testcases[180] = 76'h4202340500b3a928881;
assign testcases[181] = 76'h98035c0100d0ba3bcc4;
assign testcases[182] = 76'h7000540120814428771;
assign testcases[183] = 76'h8003660350b08629881;
assign testcases[184] = 76'h83014b0210d0b829cd8;
assign testcases[185] = 76'h8306580570d0a539984;
assign testcases[186] = 76'h8001840700824409990;
assign testcases[187] = 76'h91027244004c773dcc0;
assign testcases[188] = 76'h91037234004c773dcc1;
assign testcases[189] = 76'h92014303005a820ccb0;
assign testcases[190] = 76'h900272440095873dcc0;
assign testcases[191] = 76'hb1037104003c640dcc0;
assign testcases[192] = 76'hb1018113004d930dcc0;
assign testcases[193] = 76'hb1037104003d630dcc0;
assign testcases[194] = 76'hd0049132001e620ccc0;
assign testcases[195] = 76'hd0029122001e620ccc0;
assign testcases[196] = 76'hd002a132002e630dcc0;
assign testcases[197] = 76'hc0018114002d600ccc0;
assign testcases[198] = 76'hc1018102002e710ccc0;
assign testcases[199] = 76'h4000911410712508770;
assign testcases[200] = 76'h4000810500712408770;
assign testcases[201] = 76'h4000912300282208770;
assign testcases[202] = 76'h4000912300292028770;
assign testcases[203] = 76'h4000a10300292008770;
assign testcases[204] = 76'h4000813200291128770;
assign testcases[205] = 76'h40009122001a2008770;
assign testcases[206] = 76'h4000920500712408770;
assign testcases[207] = 76'h4000910500621308770;
assign testcases[208] = 76'h5201710200463409880;
assign testcases[209] = 76'h5000a10200292009880;
assign testcases[210] = 76'h6611810200553809980;
assign testcases[211] = 76'h61008102001b3109980;
assign testcases[212] = 76'h6401820100a17709980;
assign testcases[213] = 76'h6200710200733309980;
assign testcases[214] = 76'h6101a11300723409980;
assign testcases[215] = 76'h6101a10300394309990;
assign testcases[216] = 76'h6000b11400824409880;
assign testcases[217] = 76'h6000a11400824409880;
assign testcases[218] = 76'h640192151072382a991;
assign testcases[219] = 76'h620091060092630a990;
assign testcases[220] = 76'h7210910400734909980;
assign testcases[221] = 76'h70009102002a3309980;
assign testcases[222] = 76'h7100720500905509980;
assign testcases[223] = 76'h71007202003a5209980;
assign testcases[224] = 76'h71009102003b5309990;
assign testcases[225] = 76'h70009102002a3309980;
assign testcases[226] = 76'h6500820400724209980;
assign testcases[227] = 76'h6200820500724208981;
assign testcases[228] = 76'h6200720400723209980;
assign testcases[229] = 76'h5200910500802609880;
assign testcases[230] = 76'h5100910300654409880;
assign testcases[231] = 76'h5000811400622209880;
assign testcases[232] = 76'h5100910300654409880;
assign testcases[233] = 76'h5000811400622209880;
assign testcases[234] = 76'h5000811400622209880;
assign testcases[235] = 76'h4200910300722308880;
assign testcases[236] = 76'h41009103002a2008870;
assign testcases[237] = 76'h4200a112002a2008880;
assign testcases[238] = 76'h6001c08200292008770;
assign testcases[239] = 76'h6001c0a2001a1108770;
assign testcases[240] = 76'h6000c0d1000a1008870;
assign testcases[241] = 76'h6001c05210702408770;
assign testcases[242] = 76'h6001c04200291108770;
assign testcases[243] = 76'h5001c15400a05608770;
assign testcases[244] = 76'h5000c16300665408770;
assign testcases[245] = 76'h7503740600b19909991;
assign testcases[246] = 76'h720382040091530a990;
assign testcases[247] = 76'hd4019141003d830cdc0;
assign testcases[248] = 76'hd4018100003d820ddd0;
assign testcases[249] = 76'hd100b071002d620ccc0;
assign testcases[250] = 76'hc101a152002d620ccb0;
assign testcases[251] = 76'h7003c14500735b0aaa0;
assign testcases[252] = 76'h7103a15500825609981;
assign testcases[253] = 76'h7000919200192208770;
assign testcases[254] = 76'h7001817300293308870;
assign testcases[255] = 76'h6506070260b2a709883;
assign testcases[256] = 76'h6203080230b19709782;
assign testcases[257] = 76'h6202180040c0aa0c788;
assign testcases[258] = 76'h6403080020c0ab29882;
assign testcases[259] = 76'h6104070320925339782;
assign testcases[260] = 76'h600223040088a429980;
assign testcases[261] = 76'h600323040088a509990;
assign testcases[262] = 76'h600134050088a809990;
assign testcases[263] = 76'h600124050088a509990;
assign testcases[264] = 76'h6001240400394409880;
assign testcases[265] = 76'h70054204007aa30bcb1;
assign testcases[266] = 76'h5603720300825509980;
assign testcases[267] = 76'h5203720300814409980;
assign testcases[268] = 76'h62018102003a5209990;
assign testcases[269] = 76'h6201810300824209980;
assign testcases[270] = 76'h5706520110484108880;
assign testcases[271] = 76'h5503520000394309880;
assign testcases[272] = 76'h5101622400813a28870;
assign testcases[273] = 76'h5000420500723308870;
assign testcases[274] = 76'h5000716200713408870;
assign testcases[275] = 76'h5101520400723208870;
assign testcases[276] = 76'h5000624300713408870;
assign testcases[277] = 76'h51039123002a3408880;
assign testcases[278] = 76'h50018112002a2108870;
assign testcases[279] = 76'h4308831320a07638871;
assign testcases[280] = 76'h4204922300b19908880;
assign testcases[281] = 76'h4204650220a07508771;
assign testcases[282] = 76'h810272052067640a991;
assign testcases[283] = 76'h80007206003a5309990;
assign testcases[284] = 76'h720172020059750a990;
assign testcases[285] = 76'hb000c062002c530bbb0;
assign testcases[286] = 76'hb000d092002c430bbb0;
assign testcases[287] = 76'hb000a113003b630baa0;
assign testcases[288] = 76'hb000a103003b630aaa0;
assign testcases[289] = 76'hb000d0a1001e420bbb0;
assign testcases[290] = 76'hb000b043002c520bba0;
assign testcases[291] = 76'hb000a19400734b0aaa0;
assign testcases[292] = 76'hb000821600a17b0aaa0;
assign testcases[293] = 76'hb000a1650091590baa0;
assign testcases[294] = 76'hc000c17400a4950bba0;
assign testcases[295] = 76'hc000d1a400a4940bba0;
assign testcases[296] = 76'hc010d0e1001d400bbb0;
assign testcases[297] = 76'hc000d0f1000e410bbb0;
assign testcases[298] = 76'hc000c0c1001d410bbb0;
assign testcases[299] = 76'hc000d0a1001d410bbb0;
assign testcases[300] = 76'hb000d092001d410baa0;
assign testcases[301] = 76'hb000e0b1001d420baa0;
assign testcases[302] = 76'hb000d042001c410baa0;
assign testcases[303] = 76'hc010d072005c930baa0;
assign testcases[304] = 76'hc000e082002c410bba0;
assign testcases[305] = 76'hc010d053005c920baa0;
assign testcases[306] = 76'hc000e082002c410bba0;
assign testcases[307] = 76'h8000a062001b3109990;
assign testcases[308] = 76'ha000d0c30073320baa0;
assign testcases[309] = 76'ha000e0d1001d310baa0;
assign testcases[310] = 76'hc000c183004a550cbb0;
assign testcases[311] = 76'hc000e0a1001c420bbb0;
assign testcases[312] = 76'hc000b163003c640cbb0;
assign testcases[313] = 76'hc000d072003a540bba0;
assign testcases[314] = 76'hc000e0b2002a440bba0;
assign testcases[315] = 76'hc000c042002d510bba0;
assign testcases[316] = 76'hd010d0a2002c540bbb0;
assign testcases[317] = 76'hd000e0f1000e410bbb0;
assign testcases[318] = 76'hb010d0a2002c540bbb0;
assign testcases[319] = 76'hd000e0f1000e410bbb0;
assign testcases[320] = 76'hd000d032001d500bbb0;
assign testcases[321] = 76'hd000d082002b430bbb0;
assign testcases[322] = 76'h900092750082570aaa0;
assign testcases[323] = 76'h9000b1c20083630aaa0;
assign testcases[324] = 76'h9000b1c20083630aaa0;
assign testcases[325] = 76'h9110922500c2a90baa1;
assign testcases[326] = 76'hb000e0b30073430baa0;
assign testcases[327] = 76'hb000d0c1001d420bba0;
assign testcases[328] = 76'hc000f0e1001d410bba0;
assign testcases[329] = 76'hc000e071001d410aaa0;
assign testcases[330] = 76'hc000e0a1001d410baa0;
assign testcases[331] = 76'hc000e0a1001d410baa0;
assign testcases[332] = 76'hc000e042001d400aaa0;
assign testcases[333] = 76'hb000e0b30073430baa0;
assign testcases[334] = 76'hb000e0e20073420baa0;
assign testcases[335] = 76'hc000f0c1001d410baa0;
assign testcases[336] = 76'h9010b1230073420aaa0;
assign testcases[337] = 76'h9000b023002c410baa0;
assign testcases[338] = 76'h9000b023002c410baa0;
assign testcases[339] = 76'h8000d0f1000c2109990;
assign testcases[340] = 76'h8000d0f1000c2109990;
assign testcases[341] = 76'h8000d0e1000c2109990;
assign testcases[342] = 76'h8000d0f1000c2109990;
assign testcases[343] = 76'ha000d0830072350aa90;
assign testcases[344] = 76'ha000e072001b312aaa0;
assign testcases[345] = 76'ha000e0a1001c310aa90;
assign testcases[346] = 76'ha000e0a1001c310aa90;
assign testcases[347] = 76'ha000e022001b312aa90;
assign testcases[348] = 76'ha001e0b1001c310aaa0;
assign testcases[349] = 76'ha001e092001d310aaa0;
assign testcases[350] = 76'ha000d091001d310aaa0;
assign testcases[351] = 76'ha000e0e1000d310aaa0;
assign testcases[352] = 76'ha000e0f1000d310aa90;
assign testcases[353] = 76'ha000c043002c420aaa0;
assign testcases[354] = 76'ha000c042102b310aa90;
assign testcases[355] = 76'ha000a23430b2a82aa91;
assign testcases[356] = 76'h7000a1330057440aaa0;
assign testcases[357] = 76'h710072050081570a990;
assign testcases[358] = 76'h8002a1240073440a990;
assign testcases[359] = 76'h800191040073420aa90;
assign testcases[360] = 76'h8001b042001c320a990;
assign testcases[361] = 76'h8001c052001c310a990;
assign testcases[362] = 76'h9001c0c2002a340a990;
assign testcases[363] = 76'h9001c0e1001c310a990;
assign testcases[364] = 76'h9001c0f1001c310a990;
assign testcases[365] = 76'h9001a1430039340a990;
assign testcases[366] = 76'h9001b0b1000c310a990;
assign testcases[367] = 76'h9001b0c2002a330a990;
assign testcases[368] = 76'h8001a112001b3109990;
assign testcases[369] = 76'h9001b052203a520baa0;
assign testcases[370] = 76'h9000c042002b410baa0;
assign testcases[371] = 76'h900191031048440baa0;
assign testcases[372] = 76'h9001a1621058540baa1;
assign testcases[373] = 76'h9000c042103a420baa0;
assign testcases[374] = 76'h9001a1231048430baa0;
assign testcases[375] = 76'ha001a072103a530cbb0;
assign testcases[376] = 76'ha411925210b18c0cbb1;
assign testcases[377] = 76'ha300720100a1760cbb0;
assign testcases[378] = 76'ha101a172103a530cbb0;
assign testcases[379] = 76'ha1019132104a740cbb0;
assign testcases[380] = 76'ha301820110a1760bbb0;
assign testcases[381] = 76'h7712620100c2b429ba4;
assign testcases[382] = 76'h7611530100c2b42aca4;
assign testcases[383] = 76'h72107101006b910ab92;
assign testcases[384] = 76'h81008102002b4109990;
assign testcases[385] = 76'h7612530610c2aa3fca9;
assign testcases[386] = 76'h731153000097a32fde6;
assign testcases[387] = 76'h720152030096a70fcb8;
assign testcases[388] = 76'h7100620400915338991;
assign testcases[389] = 76'h7211530400c1a66fbab;
assign testcases[390] = 76'h7411530300c1a45aba3;
assign testcases[391] = 76'hb001a153003a542bba0;
assign testcases[392] = 76'hb000c092001d410baa0;
assign testcases[393] = 76'hb001720400a3942bbb0;
assign testcases[394] = 76'hb001912400a3942bba0;
assign testcases[395] = 76'hb001b163003a542bba0;
assign testcases[396] = 76'hb001812400a3952bba0;
assign testcases[397] = 76'hc000b042002d610ccc0;
assign testcases[398] = 76'hc000b042001e600ccc0;
assign testcases[399] = 76'hd100732420d0a70ccc1;
assign testcases[400] = 76'hd00091b1001f600ddc0;
assign testcases[401] = 76'hd000723210c2a40ccc0;
assign testcases[402] = 76'hd00081c1000f600ccc0;
assign testcases[403] = 76'hd00071c1000f600ccc0;
assign testcases[404] = 76'hd000d28230d0b70cbb2;
assign testcases[405] = 76'hd000c38130d0b90cbb3;
assign testcases[406] = 76'hd000e092001e510ccb0;
assign testcases[407] = 76'hd000e052001e510ccb0;
assign testcases[408] = 76'hd000e082103b510ccb0;
assign testcases[409] = 76'hd000e092001e500ccb0;
assign testcases[410] = 76'hc001c0320074410bba0;
assign testcases[411] = 76'hc001d032101d400aba0;
assign testcases[412] = 76'hc000a022001e400bbb0;
assign testcases[413] = 76'hc000b0230074410bbb0;
assign testcases[414] = 76'h9101a11300a3930aa90;
assign testcases[415] = 76'h90009102002c4209a90;
assign testcases[416] = 76'h9100b112003c610aaa0;
assign testcases[417] = 76'h9101c082006cb30aaa0;
assign testcases[418] = 76'h9000d0c1001c410aaa0;
assign testcases[419] = 76'h9101b122007bb40baa0;
assign testcases[420] = 76'h9100c081006cb30aaa0;
assign testcases[421] = 76'hb003b124003a540bba0;
assign testcases[422] = 76'hb001b1540073562bba0;
assign testcases[423] = 76'hb001b103002c422aaa0;
assign testcases[424] = 76'hb001b114002c542bba0;
assign testcases[425] = 76'hf0019113002d622ddc0;
assign testcases[426] = 76'hf00391160088a30ddc0;
assign testcases[427] = 76'h4902630200835429991;
assign testcases[428] = 76'h450163020098b629980;
assign testcases[429] = 76'h4601630200c3b729980;
assign testcases[430] = 76'h4701620200834629990;
assign testcases[431] = 76'h660062040057540a990;
assign testcases[432] = 76'h6500530400b3a328981;
assign testcases[433] = 76'h63007202003a530a990;
assign testcases[434] = 76'hd005b34370d0b75cbc3;
assign testcases[435] = 76'hd002a23120b0770cbb2;
assign testcases[436] = 76'hd003b25140d0ba3cbc2;
assign testcases[437] = 76'hd004a33340d0b72cbb2;
assign testcases[438] = 76'hd004a63940d0bbdcbc3;
assign testcases[439] = 76'hd003961740d0babcbb4;
assign testcases[440] = 76'hb101932520a06b5baa1;
assign testcases[441] = 76'hb101932320a06d5baa1;
assign testcases[442] = 76'hb000a11310a1630bbb1;
assign testcases[443] = 76'hb000a012001d500bbb0;
assign testcases[444] = 76'hb000a112002d610bbb0;
assign testcases[445] = 76'hb000c072001d410aaa0;
assign testcases[446] = 76'hb000c072001d410aaa0;
assign testcases[447] = 76'hb000c072001d410aaa0;
assign testcases[448] = 76'h9300a1220083640aaa0;
assign testcases[449] = 76'h9100a1330083640aa90;
assign testcases[450] = 76'h9000a1330039440aa90;
assign testcases[451] = 76'h9300a1110083640aaa0;
assign testcases[452] = 76'h6603740600b19909991;
assign testcases[453] = 76'h80019133002b310a990;
assign testcases[454] = 76'h8001a133002b320a990;
assign testcases[455] = 76'h80019123002b320a990;
assign testcases[456] = 76'h7413550610905209991;
assign testcases[457] = 76'ha401640500a3972cbb1;
assign testcases[458] = 76'ha20072050093710cbb0;
assign testcases[459] = 76'ha20171130093630aba0;
assign testcases[460] = 76'h4201b02200383208770;
assign testcases[461] = 76'h4000c04200192208760;
assign testcases[462] = 76'h4201910300383108870;
assign testcases[463] = 76'h4401831400a17e27881;
assign testcases[464] = 76'h4101911300836607871;
assign testcases[465] = 76'hb001e14310b4b40bba0;
assign testcases[466] = 76'hb001f052003c720baa0;
assign testcases[467] = 76'hb001f052003c720baa0;
assign testcases[468] = 76'hb001f062003c720baa0;
assign testcases[469] = 76'hd000f052003c620ccb0;
assign testcases[470] = 76'hd000f052002c520cbb0;
assign testcases[471] = 76'hd000f072001e500ccb0;
assign testcases[472] = 76'hd001f032004c720cbb0;
assign testcases[473] = 76'hd000f043004b710bcb0;
assign testcases[474] = 76'hd000f062002d500bbb0;
assign testcases[475] = 76'hd000f072001d500bbb0;
assign testcases[476] = 76'hc001b1131083512bba0;
assign testcases[477] = 76'hc000c022002c510bbb0;
assign testcases[478] = 76'hc001a1121049512bba0;
assign testcases[479] = 76'hc000a1021049512bbb0;
assign testcases[480] = 76'ha001a16400b4b80aaa0;
assign testcases[481] = 76'ha000b1720075540aaa0;
assign testcases[482] = 76'ha1009113005b962bba0;
assign testcases[483] = 76'ha100921300b1752cba1;
assign testcases[484] = 76'hb001a1350074592baa0;
assign testcases[485] = 76'hb000b032001d420baa0;
assign testcases[486] = 76'h6600520210a28509a82;
assign testcases[487] = 76'h6400520100b28509a92;
assign testcases[488] = 76'h6200430210847409982;
assign testcases[489] = 76'h6600520100a28509a92;
assign testcases[490] = 76'h4821550400b1790dbc4;
assign testcases[491] = 76'h4610460300d0a80dbc5;
assign testcases[492] = 76'h4621540000c0ac0dbc3;
assign testcases[493] = 76'h4421540300b0850dcc2;
assign testcases[494] = 76'h6711550200a27c29aa2;
assign testcases[495] = 76'h6411630200a27529a93;
assign testcases[496] = 76'h7a31450300b0790cbb2;
assign testcases[497] = 76'h7621540100c0870cbb1;
assign testcases[498] = 76'h7830460400b07b0cbc1;
assign testcases[499] = 76'h7721540200c0890cbb2;
assign testcases[500] = 76'h7a11480200b07a2bab2;
assign testcases[501] = 76'h7701470200c0992bab1;
assign testcases[502] = 76'h7603540600a1750cbb2;
assign testcases[503] = 76'h7403540500a0740cbb2;
assign testcases[504] = 76'h7402620400b18609a91;
assign testcases[505] = 76'h7202620400b18709a91;
assign testcases[506] = 76'hf6018102003fa00ded0;
assign testcases[507] = 76'hf4018102003fa10ded0;
assign testcases[508] = 76'hf5018102003fa10ded0;
assign testcases[509] = 76'hf3018101003fa20ded1;
assign testcases[510] = 76'he4028102006b933ddd0;
assign testcases[511] = 76'he4017101004e922ded1;
assign testcases[512] = 76'he1019103003d710ddc0;
assign testcases[513] = 76'he1009102002f812ddc0;
assign testcases[514] = 76'h7614720200835429aa1;
assign testcases[515] = 76'h7212710200835309a91;
assign testcases[516] = 76'h7302620100948309a91;
assign testcases[517] = 76'h7412720100a3830caa1;
assign testcases[518] = 76'h6413630300b2a809981;
assign testcases[519] = 76'h6312630200d0a809981;
assign testcases[520] = 76'h6101621400824309880;
assign testcases[521] = 76'h60006213002a3129880;
assign testcases[522] = 76'hf6116204004fa40fff1;
assign testcases[523] = 76'hf4116100004fa20fff1;
assign testcases[524] = 76'hf4116200003fa10fff1;
assign testcases[525] = 76'hf3006201004fa20fff1;
assign testcases[526] = 76'hbb21540110d0bb0fde3;
assign testcases[527] = 76'hb6116300005b970fef1;
assign testcases[528] = 76'hb41162000079920fff1;
assign testcases[529] = 76'hb410450000d1b90ecc2;
assign testcases[530] = 76'hb410470110d0b90dcc3;
assign testcases[531] = 76'hb611630000b3a40fff1;
assign testcases[532] = 76'h9200a1440083670aaa0;
assign testcases[533] = 76'h9000a1440083630aaa0;
assign testcases[534] = 76'h9000b1620083630aaa0;
assign testcases[535] = 76'h910092350094772aaa0;
assign testcases[536] = 76'h910091420094740aaa0;
assign testcases[537] = 76'hb000b1550083640baa0;
assign testcases[538] = 76'hb000c1540083640baa0;
assign testcases[539] = 76'hb000b14300a1640aaa0;
assign testcases[540] = 76'hc40181030084640ccc0;
assign testcases[541] = 76'hc1009102002e600ccc0;
assign testcases[542] = 76'ha10191050091660bba0;
assign testcases[543] = 76'ha00191050073540aba0;
assign testcases[544] = 76'hc000c052102b440bba0;
assign testcases[545] = 76'hc001c072001d410bba0;
assign testcases[546] = 76'hc000b043003b440baa0;
assign testcases[547] = 76'h9012a1521057440bba0;
assign testcases[548] = 76'ha003a133002c410baa0;
assign testcases[549] = 76'ha001a042001c410baa0;
assign testcases[550] = 76'ha002a142002b410baa0;
assign testcases[551] = 76'h97055d0900d0b45bbb4;
assign testcases[552] = 76'h97025b0200d0ba3bdc4;
assign testcases[553] = 76'ha2075b0940b0792baa3;
assign testcases[554] = 76'ha003590740b0882a9a2;
assign testcases[555] = 76'ha2036c0b00d0b72bbb3;
assign testcases[556] = 76'ha104680730b0840aaa1;
assign testcases[557] = 76'h7202660920d0a539992;
assign testcases[558] = 76'h7202550320d0a639982;
assign testcases[559] = 76'h7101560420d0a728983;
assign testcases[560] = 76'h7000540120814428771;
assign testcases[561] = 76'h7108560530c1a829882;
assign testcases[562] = 76'h7004740430a06729771;
assign testcases[563] = 76'h7105470520c0a908974;
assign testcases[564] = 76'h7103380610c1a828985;
assign testcases[565] = 76'h7504760340b08829991;
assign testcases[566] = 76'h7302750140d0ba29881;
assign testcases[567] = 76'h7303841220c0a709991;
assign testcases[568] = 76'h7303650140d0bb39881;
assign testcases[569] = 76'h7506580560d0a539984;
assign testcases[570] = 76'h7103660640b08509881;
assign testcases[571] = 76'h7403580630d0b629a95;
assign testcases[572] = 76'h7404580640d0a639a95;
assign testcases[573] = 76'h7303590810d0b629b96;
assign testcases[574] = 76'h73015b0510d0b639cd8;
assign testcases[575] = 76'h7003660540b08429781;
assign testcases[576] = 76'h7103660540b08609881;
assign testcases[577] = 76'h9200c10510b1840aa90;
assign testcases[578] = 76'h4203620300687508972;
assign testcases[579] = 76'h4001710400292208770;
assign testcases[580] = 76'h4101520300292108880;
assign testcases[581] = 76'h4203620300687408871;
assign testcases[582] = 76'h4101620300697408972;
assign testcases[583] = 76'h4203620300697608972;
assign testcases[584] = 76'h4102620410a17907761;
assign testcases[585] = 76'h4001720310383307660;
assign testcases[586] = 76'h4001620400282108760;
assign testcases[587] = 76'h4213530400a27507872;
assign testcases[588] = 76'h4001630500586507760;
assign testcases[589] = 76'h4001630500586407760;
assign testcases[590] = 76'h4213540300b29608983;
assign testcases[591] = 76'h410253050077742da94;
assign testcases[592] = 76'h420253010084760da94;
assign testcases[593] = 76'h4202530400847407973;
assign testcases[594] = 76'hc103e113003d720bcb0;
assign testcases[595] = 76'hc003e013002d510bbb0;
assign testcases[596] = 76'hc002f013001e500bbb0;
assign testcases[597] = 76'hc002e113003d710bbb0;
assign testcases[598] = 76'hc003e113003d710bbb0;
assign testcases[599] = 76'hc001d103003d710bbb0;
assign testcases[600] = 76'hb401d1031085740ccb0;
assign testcases[601] = 76'hb101e104005b820ccb0;
assign testcases[602] = 76'hb401d1011085730ccb0;
assign testcases[603] = 76'hb401d1021095830ccc0;
assign testcases[604] = 76'hb200c2030093740bbb0;
assign testcases[605] = 76'hc602d103007aa20ccc1;
assign testcases[606] = 76'hc201c103006aa10ccc1;
assign testcases[607] = 76'hc402d103007aa20cdc1;
assign testcases[608] = 76'hb40253060093742bbb1;
assign testcases[609] = 76'hb301530400a1722bbb1;
assign testcases[610] = 76'hb101540800a1752bbb1;
assign testcases[611] = 76'hb30144070093742bbb1;
assign testcases[612] = 76'hb101630300c1a82bbb0;
assign testcases[613] = 76'hc701640900b0860ccb1;
assign testcases[614] = 76'hc501640800b0740cbb1;
assign testcases[615] = 76'hc401640800c0870ccc1;
assign testcases[616] = 76'hc811620000a3930cdd1;
assign testcases[617] = 76'hb001461c0090510aaa1;
assign testcases[618] = 76'hb00062230081420baa0;
assign testcases[619] = 76'hb603720300c0840bcb1;
assign testcases[620] = 76'hb602720100c0940ccc1;
assign testcases[621] = 76'hb0017113002d620bba0;
assign testcases[622] = 76'h861357090091540a9a2;
assign testcases[623] = 76'h8401650600a1630a991;
assign testcases[624] = 76'h7512760900a06209991;
assign testcases[625] = 76'h7412750900a06209a91;
assign testcases[626] = 76'h8300550510a0690aaa2;
assign testcases[627] = 76'h4201732610c19808771;
assign testcases[628] = 76'h40018152002a2008770;
assign testcases[629] = 76'h8a03760030a1740bbb2;
assign testcases[630] = 76'h8902850000b0740dbb2;
assign testcases[631] = 76'hb000822700a3980cbb0;
assign testcases[632] = 76'hb00071240084642cbb0;
assign testcases[633] = 76'hb000b112001e510ccb0;
assign testcases[634] = 76'hb200821410b4b70bbb0;
assign testcases[635] = 76'hb000a1130094720bbb0;
assign testcases[636] = 76'hb00091030058630bbb0;
assign testcases[637] = 76'hb20073040094850bba0;
assign testcases[638] = 76'h9300720400a3960baa0;
assign testcases[639] = 76'h9200620400a3940baa0;
assign testcases[640] = 76'h900062050073540baa0;
assign testcases[641] = 76'h900062060083530baa0;
assign testcases[642] = 76'h9600650600c0948baa1;
assign testcases[643] = 76'h9400730200d0bb0bba0;
assign testcases[644] = 76'h5001d0d200292308770;
assign testcases[645] = 76'h5000e0f1001a1108770;
assign testcases[646] = 76'h5001a10300452408770;
assign testcases[647] = 76'h5001d0b200452308770;
assign testcases[648] = 76'h5001d0a200452308770;
assign testcases[649] = 76'h5000c0c200271108770;
assign testcases[650] = 76'h5000d0f1001a1208770;
assign testcases[651] = 76'h5000d0f1001a1208770;
assign testcases[652] = 76'h5000c09200371008770;
assign testcases[653] = 76'h5000c0c100191208770;
assign testcases[654] = 76'h5000d0e100191108770;
assign testcases[655] = 76'h7204232300825609980;
assign testcases[656] = 76'h7203231300a28809990;
assign testcases[657] = 76'h71032322003a4209980;
assign testcases[658] = 76'h71023222003a5109990;
assign testcases[659] = 76'h71022322003a4109980;
assign testcases[660] = 76'h71022322003a4209980;
assign testcases[661] = 76'h70012e0054d0a934426;
assign testcases[662] = 76'h9003a32318c1a82a894;
assign testcases[663] = 76'h9003a32318c1aa2a894;
assign testcases[664] = 76'h9001a21204a3992a894;
assign testcases[665] = 76'h9002a22304a39b2a893;
assign testcases[666] = 76'h9001b123002a410aaa0;
assign testcases[667] = 76'h9001b022002c430aaa0;
assign testcases[668] = 76'h9002a23214c1a73a993;
assign testcases[669] = 76'ha101921330b19b3baa3;
assign testcases[670] = 76'ha101922330c1a73b9a4;
assign testcases[671] = 76'ha00071031058552caa1;
assign testcases[672] = 76'ha101b122003b510bbb0;
assign testcases[673] = 76'ha901a30100c0940fdd2;
assign testcases[674] = 76'ha601a30300c0940fde2;
assign testcases[675] = 76'ha600930000c0930bdd2;
assign testcases[676] = 76'ha400a200005a810fde2;
assign testcases[677] = 76'ha600930000c0930fdd2;
assign testcases[678] = 76'ha400a20100b2940fde2;
assign testcases[679] = 76'hb10382080091670baa0;
assign testcases[680] = 76'hb1019103004a730bba0;
assign testcases[681] = 76'ha203560d00a2883bba1;
assign testcases[682] = 76'h8051560028d1b832206;
assign testcases[683] = 76'h8041550018a16422205;
assign testcases[684] = 76'h825633052066510a991;
assign testcases[685] = 76'h824433042083520a991;
assign testcases[686] = 76'h8001430500393109990;
assign testcases[687] = 76'h823333042066520a991;
assign testcases[688] = 76'h824333031083520a991;
assign testcases[689] = 76'h83e325054492760a895;
assign testcases[690] = 76'h8051160714927407763;
assign testcases[691] = 76'h828134042093762a992;
assign testcases[692] = 76'h8382340430b0850a894;
assign testcases[693] = 76'h83f4440344a18629882;
assign testcases[694] = 76'h8292530220835609991;
assign testcases[695] = 76'h8193340234915409782;
assign testcases[696] = 76'h8282430310835409991;
assign testcases[697] = 76'h71d3440348a16c09676;
assign testcases[698] = 76'h7061550124b18922449;
assign testcases[699] = 76'h7192340344c1ae09882;
assign testcases[700] = 76'h709245023cc19c09578;
assign testcases[701] = 76'h7051a40414b19a09783;
assign testcases[702] = 76'h7030f00204473306873;
assign testcases[703] = 76'h7030f00204473306772;
assign testcases[704] = 76'h7020f00004282106761;
assign testcases[705] = 76'h8006a1a300b3b729980;
assign testcases[706] = 76'h8004b0e1001b2109980;
assign testcases[707] = 76'h71069113002a3209980;
assign testcases[708] = 76'h70039122002b3109980;
assign testcases[709] = 76'h60049152002a3209880;
assign testcases[710] = 76'h60019172002a3209880;
assign testcases[711] = 76'h6203640820b07729881;
assign testcases[712] = 76'h6202640700904409881;
assign testcases[713] = 76'h4201731600905709881;
assign testcases[714] = 76'h84059133004a5209a90;
assign testcases[715] = 76'h83039103004a520aaa0;
assign testcases[716] = 76'h8103a142003a5209980;
assign testcases[717] = 76'h8001b072002a3209980;
assign testcases[718] = 76'h81018104003a522a990;
assign testcases[719] = 76'h7003b092002a3109880;
assign testcases[720] = 76'h7001b0d1000b2109880;
assign testcases[721] = 76'hb010b082002c520bba0;
assign testcases[722] = 76'hb000c092001e510bba0;
assign testcases[723] = 76'hb0109114004a540bba0;
assign testcases[724] = 76'h74129102003a540aa90;
assign testcases[725] = 76'h72029102003a530aa90;
assign testcases[726] = 76'h700191030057530aa90;
assign testcases[727] = 76'h72019101003a5009a91;
assign testcases[728] = 76'h4203811200814208870;
assign testcases[729] = 76'h4202811200814208871;
assign testcases[730] = 76'h40019113001a2108770;
assign testcases[731] = 76'h42017103004a520caa2;
assign testcases[732] = 76'h41028112003a4308870;
assign testcases[733] = 76'h56166303006a982bbb1;
assign testcases[734] = 76'h7411720200a4950baa1;
assign testcases[735] = 76'h76136302006a992bbb1;
assign testcases[736] = 76'h74146303006a982bbb1;
assign testcases[737] = 76'h5603640700813608881;
assign testcases[738] = 76'h5401630500803529881;
assign testcases[739] = 76'h4401651800916428771;
assign testcases[740] = 76'h4400640600916409881;
assign testcases[741] = 76'ha20191120092620bba0;
assign testcases[742] = 76'ha101a012001d510bba0;
assign testcases[743] = 76'hb1033701b0c0973a893;
assign testcases[744] = 76'hb0010a0050b08c55665;
assign testcases[745] = 76'hb103280190d0ab2a894;
assign testcases[746] = 76'hb103460180d0a70a992;
assign testcases[747] = 76'hb103370180d0a60a893;
assign testcases[748] = 76'h8000e072001b3209990;
assign testcases[749] = 76'h8000f092001c3209990;
assign testcases[750] = 76'h8000f0b1001c3109990;
assign testcases[751] = 76'h8000e072001b3209990;
assign testcases[752] = 76'h71009162005b8409980;
assign testcases[753] = 76'h70009162001b3209980;
assign testcases[754] = 76'h7000a062002b3109980;
assign testcases[755] = 76'h7000a072002b3209980;
assign testcases[756] = 76'h7000721700803309880;
assign testcases[757] = 76'h7000822400622109880;
assign testcases[758] = 76'h7200a10300b29629980;
assign testcases[759] = 76'h7000c003002b3009980;
assign testcases[760] = 76'h7200a0120069840aa90;
assign testcases[761] = 76'h7200a012002a420a990;
assign testcases[762] = 76'h7000c022002b400a990;
assign testcases[763] = 76'h7200a24600a29f09990;
assign testcases[764] = 76'ha000c0830073420aaa0;
assign testcases[765] = 76'ha000e0b1001c310aaa0;
assign testcases[766] = 76'ha000a052001c410baa0;
assign testcases[767] = 76'h9000c0c10072320a990;
assign testcases[768] = 76'h9000c0d1001c310a990;
assign testcases[769] = 76'h8000f0f0000c2109990;
assign testcases[770] = 76'h8000f0f0000c2109990;
assign testcases[771] = 76'h7000e0f110282509880;
assign testcases[772] = 76'h7000d07110586509880;
assign testcases[773] = 76'h7000e0f1000b2109880;
assign testcases[774] = 76'h7000d0c110586509880;
assign testcases[775] = 76'h9001e072002b520aa90;
assign testcases[776] = 76'h9001d062002b420aa90;
assign testcases[777] = 76'h9001d062002b420aa90;
assign testcases[778] = 76'h9001d052002b420aa90;
assign testcases[779] = 76'h7000d062002b3109980;
assign testcases[780] = 76'h7000d072002b3109880;
assign testcases[781] = 76'h7000e062001b3209990;
assign testcases[782] = 76'h7000d082002b3109880;
assign testcases[783] = 76'h8000c043005b9409990;
assign testcases[784] = 76'h8000d043003a3209990;
assign testcases[785] = 76'h3100911400712508770;
assign testcases[786] = 76'h3000812400712408770;
assign testcases[787] = 76'h5200910500802609880;
assign testcases[788] = 76'h5200911500722608880;
assign testcases[789] = 76'h5100910200654408880;
assign testcases[790] = 76'h5100821500712609880;
assign testcases[791] = 76'h5100821500712609880;
assign testcases[792] = 76'hc10c91635066640bbb0;
assign testcases[793] = 76'hc10991635066630cbb1;
assign testcases[794] = 76'hc10882635075630cbb1;
assign testcases[795] = 76'hc004b052001d520bbb0;
assign testcases[796] = 76'hc003c062001d510bbb0;
assign testcases[797] = 76'hc003b072001d510bbb0;
assign testcases[798] = 76'hc003b072001d510bbb0;
assign testcases[799] = 76'hc004b082002c530cbb0;
assign testcases[800] = 76'hc003c0a1001e500cbb0;
assign testcases[801] = 76'hc005b072102c640cbb0;
assign testcases[802] = 76'hc003b062002c610bbb0;
assign testcases[803] = 76'hc00234325075640baa2;
assign testcases[804] = 76'hc10334245075630baa1;
assign testcases[805] = 76'hc0018153004a630dcc0;
assign testcases[806] = 76'hc0019163002d622dcc0;
assign testcases[807] = 76'hc0019163002d622dcc0;
assign testcases[808] = 76'hc20462625085722cbc1;
assign testcases[809] = 76'hc001a092004a640ccc0;
assign testcases[810] = 76'hc00191831066642ccc0;
assign testcases[811] = 76'hc20353523076723dcc1;
assign testcases[812] = 76'hc20362622076725dcc1;
assign testcases[813] = 76'hc20343424085712dbc2;
assign testcases[814] = 76'hc10133022084740bbb2;
assign testcases[815] = 76'hc00133322074640bbb1;
assign testcases[816] = 76'hc10133322074640bbb1;
assign testcases[817] = 76'he001a0a3003b620dcc0;
assign testcases[818] = 76'he001a193003b620dcc0;
assign testcases[819] = 76'he002a0b2003c632dcc0;
assign testcases[820] = 76'he001a0a2003c632dcc0;
assign testcases[821] = 76'he002b0c1001f610dcc0;
assign testcases[822] = 76'he002a0b1001f610dcc0;
assign testcases[823] = 76'he002a0c2002c640dcc0;
assign testcases[824] = 76'he001a0d2003b640dcc0;
assign testcases[825] = 76'he003b0a2002d500ccc0;
assign testcases[826] = 76'he003a1821059645ccc0;
assign testcases[827] = 76'he00291821067645ccc0;
assign testcases[828] = 76'he002a1b3003b632dcc0;
assign testcases[829] = 76'he003a1a21059633ccc0;
assign testcases[830] = 76'he003a1921059645ccc0;
assign testcases[831] = 76'he001a1b11057545ccc0;
assign testcases[832] = 76'he00391721057533ccc0;
assign testcases[833] = 76'he001a183003b640dcc0;
assign testcases[834] = 76'h740225015093762caa3;
assign testcases[835] = 76'h7201170150a1752a892;
assign testcases[836] = 76'h710126044084722b9a2;
assign testcases[837] = 76'h740135024084722caa3;
assign testcases[838] = 76'h900371a20039430aa90;
assign testcases[839] = 76'h900371b20039430aa90;
assign testcases[840] = 76'h900171920039440aa90;
assign testcases[841] = 76'h900161820039430aaa0;
assign testcases[842] = 76'h900361820039420aaa0;
assign testcases[843] = 76'h900271b2001c410aaa0;
assign testcases[844] = 76'h90027192001c410aaa0;
assign testcases[845] = 76'h910261230048440aaa0;
assign testcases[846] = 76'h910361230048440aaa0;
assign testcases[847] = 76'h910361130048440aaa0;
assign testcases[848] = 76'h910361130048540aaa0;
assign testcases[849] = 76'h910361130048540aaa0;
assign testcases[850] = 76'h91027123002c500aaa0;
assign testcases[851] = 76'h91037122002c500bba0;
assign testcases[852] = 76'h90016123002c420aaa0;
assign testcases[853] = 76'h90016172002c420aa90;
assign testcases[854] = 76'h900171a2001c310aaa0;
assign testcases[855] = 76'hb0027143002c510baa0;
assign testcases[856] = 76'hb0017113002c510baa0;
assign testcases[857] = 76'hb0037104003b510bba0;
assign testcases[858] = 76'hb0036104003b500bba0;
assign testcases[859] = 76'hb0016204003b500bbb0;
assign testcases[860] = 76'hb1026204003b510bbb0;
assign testcases[861] = 76'hb1027152002c510bbb0;
assign testcases[862] = 76'hb10252240083640bba0;
assign testcases[863] = 76'hb1037172002c530bba0;
assign testcases[864] = 76'hb1017133002c500bbb0;
assign testcases[865] = 76'hb1016204003b510bbb0;
assign testcases[866] = 76'hb0018152001d510bbb0;
assign testcases[867] = 76'hb1037172002c530bba0;
assign testcases[868] = 76'hb1037172003a540bba0;
assign testcases[869] = 76'h95046141003a520aaa0;
assign testcases[870] = 76'h94036141003a522aaa0;
assign testcases[871] = 76'h92026131003a520aaa0;
assign testcases[872] = 76'h92036141003a530aaa0;
assign testcases[873] = 76'h91027131002c510aaa0;
assign testcases[874] = 76'h91027122002b420aaa0;
assign testcases[875] = 76'h91036113003a430aaa0;
assign testcases[876] = 76'h91036113003a430aaa0;
assign testcases[877] = 76'h91036113003a420aa90;
assign testcases[878] = 76'h910362140048410aa90;
assign testcases[879] = 76'h91035204003a420aa90;
assign testcases[880] = 76'h910252040048420aa90;
assign testcases[881] = 76'h900362040039430aa90;
assign testcases[882] = 76'h91035203002b420aa90;
assign testcases[883] = 76'h91035223003b530aa90;
assign testcases[884] = 76'h91026152003b540aa90;
assign testcases[885] = 76'h90017182001c310aaa0;
assign testcases[886] = 76'h91037181001c420aaa0;
assign testcases[887] = 76'h90038142001c410baa0;
assign testcases[888] = 76'h90029152001d410baa0;
assign testcases[889] = 76'h91027181001d410aaa0;
assign testcases[890] = 76'h91037172001d410aaa0;
assign testcases[891] = 76'h90038152001d410baa0;
assign testcases[892] = 76'h91037172002c430aaa0;
assign testcases[893] = 76'hb0036113002c510bbb0;
assign testcases[894] = 76'hb0045103002c500bba0;
assign testcases[895] = 76'hb0045214002c500bbb0;
assign testcases[896] = 76'hb1055203003b500bbb0;
assign testcases[897] = 76'hb0034204003b510bbb0;
assign testcases[898] = 76'hb1034204004b600bbb0;
assign testcases[899] = 76'hb1024204005a740bbb0;
assign testcases[900] = 76'hb1024306005a730bbb1;
assign testcases[901] = 76'hb10433072077732bbb1;
assign testcases[902] = 76'hb00324072077733baa1;
assign testcases[903] = 76'hc00533271076752bbb0;
assign testcases[904] = 76'hc00543162076640bba0;
assign testcases[905] = 76'hc00342013057530baa0;
assign testcases[906] = 76'hc20342023058623bbb0;
assign testcases[907] = 76'hc20343022067622bbb0;
assign testcases[908] = 76'hc6063302006a962ccb0;
assign testcases[909] = 76'hc2033303005b940ccc0;
assign testcases[910] = 76'hc100180550d0b72baa2;
assign testcases[911] = 76'hc20135045084772cbb2;
assign testcases[912] = 76'hc2033305105a740ccb0;
assign testcases[913] = 76'h5001612300281108770;
assign testcases[914] = 76'h5001510300371208770;
assign testcases[915] = 76'h5101420300473328770;
assign testcases[916] = 76'h5101330104553128771;
assign testcases[917] = 76'h5002421204553438661;
assign testcases[918] = 76'h5001522210451208661;
assign testcases[919] = 76'h5002612300281108760;
assign testcases[920] = 76'h5003512300292208870;
assign testcases[921] = 76'h5003421320372208770;
assign testcases[922] = 76'h5101420304553228771;
assign testcases[923] = 76'h5101430300473228770;
assign testcases[924] = 76'h5202420220564209881;
assign testcases[925] = 76'h5103241320655308771;
assign testcases[926] = 76'h5002331410563408770;
assign testcases[927] = 76'h5103330230665208771;
assign testcases[928] = 76'h5103330330463308771;
assign testcases[929] = 76'h5202420220564209881;
assign testcases[930] = 76'h5203520300574329980;
assign testcases[931] = 76'h5004430430462108770;
assign testcases[932] = 76'h5005520400292108870;
assign testcases[933] = 76'h5103331320665308771;
assign testcases[934] = 76'h610334052090430a881;
assign testcases[935] = 76'h610342031047332a980;
assign testcases[936] = 76'h6004420400393109980;
assign testcases[937] = 76'h6005520500393109980;
assign testcases[938] = 76'h6005520500393109980;
assign testcases[939] = 76'h900392622084645a991;
assign testcases[940] = 76'h9001c0b2002b410aaa0;
assign testcases[941] = 76'h9103a183003b580aa90;
assign testcases[942] = 76'h92039133004a560aa90;
assign testcases[943] = 76'h92019113004a610bbb0;
assign testcases[944] = 76'h9101350048a06538673;
assign testcases[945] = 76'h9200723120a0655bab2;
assign testcases[946] = 76'hb00343153074540baa1;
assign testcases[947] = 76'hb20543053074542baa1;
assign testcases[948] = 76'hb30171040049543bbb0;
assign testcases[949] = 76'hb20161030058560bbb0;
assign testcases[950] = 76'hb20452060066542bbb0;
assign testcases[951] = 76'hb00142080066520bba1;
assign testcases[952] = 76'h960452023082540baa1;
assign testcases[953] = 76'h930252034082520a991;
assign testcases[954] = 76'h900552044083530a991;
assign testcases[955] = 76'h900543064092660a991;
assign testcases[956] = 76'h9005430460836409991;
assign testcases[957] = 76'h9003430350734429991;
assign testcases[958] = 76'h900342053082440a991;
assign testcases[959] = 76'h800426076092560a893;
assign testcases[960] = 76'h800326066092560a784;
assign testcases[961] = 76'h800453193082560a991;
assign testcases[962] = 76'h810143149082450a892;
assign testcases[963] = 76'h800153156073440a891;
assign testcases[964] = 76'h830334064082442a992;
assign testcases[965] = 76'h810233053081443a992;
assign testcases[966] = 76'h820244071082483a991;
assign testcases[967] = 76'h820134061082483a991;
assign testcases[968] = 76'h800352091082582a991;
assign testcases[969] = 76'h800362190065573a990;
assign testcases[970] = 76'h800171261065320a990;
assign testcases[971] = 76'h7004441190916629784;
assign testcases[972] = 76'h700435117091662a785;
assign testcases[973] = 76'h7003441160815329784;
assign testcases[974] = 76'h7001621140633409782;
assign testcases[975] = 76'h700345225091652a895;
assign testcases[976] = 76'h710362214090450a992;
assign testcases[977] = 76'h700362223090460a993;
assign testcases[978] = 76'h7203440174b0860a895;
assign testcases[979] = 76'h7201540034b0852a8a5;
assign testcases[980] = 76'h720263014081440a9a4;
assign testcases[981] = 76'h720262012074420a9a1;
assign testcases[982] = 76'h70034204003a4009980;
assign testcases[983] = 76'h70024204003a3009980;
assign testcases[984] = 76'h71014204002b400a990;
assign testcases[985] = 76'h74033302004a510aa90;
assign testcases[986] = 76'h73033302004a520aa90;
assign testcases[987] = 76'h77043301004a770aba0;
assign testcases[988] = 76'h750343010085770aba1;
assign testcases[989] = 76'h77032302004b730bbb0;
assign testcases[990] = 76'h740133020085850aaa1;
assign testcases[991] = 76'h740133020075640aa91;
assign testcases[992] = 76'h76033303004a760bba0;
assign testcases[993] = 76'h760333010085760aba0;
assign testcases[994] = 76'h7201320200575309980;
assign testcases[995] = 76'h71003202002b4109980;
assign testcases[996] = 76'h7403330410586409981;
assign testcases[997] = 76'h74032304004a5109a91;
assign testcases[998] = 76'h7402330400495109a91;
assign testcases[999] = 76'h780523000059640baa0;


  
  localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
  wire [$clog2(CLASS_CNT)-1:0] prediction;

  // Instantiate module under test
 cardio_tnn1_tnnseq #(
 ) dut (
    .data(data),
    .clk(clk),
    .rst(rst),
    .prediction(prediction)
  );
  
  always #halfT clk <= ~clk;

  integer i;
  initial begin
    $write("["); //" 
    for(i=0;i<TEST_CNT;i=i+1)
        runtestcase(i);
    $display("]");
    $finish;
  end

  task runtestcase(input integer i); begin
    data <= testcases[i];
    rst <= 1;
    clk <= 0;
    #period
    rst <= 0;
    #period
    #((FEAT_CNT+HIDDEN_CNT-1)*period)
    $write("%d, ",prediction);
  end
  endtask

endmodule
