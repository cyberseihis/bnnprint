












module pendigits_bs #(

parameter N = 16,
parameter M = 40,
parameter B = 4,
parameter C = 10,
parameter Ts = 5


  ) (
  input clk,
  input rst,
  input [N*B-1:0] data,
  output [$clog2(C)-1:0] klass
  );

  localparam Weights0 = 640'b0001000011111110110111111111000000010111110001101101011010000000001100111000010100010010101011010001010101000100000101000101101111100011110100100110101011001010011010110011010011110001111010111111001000111101100011110001000111010100011100011011110000011001011010010000101111111011001110000000100100101101110001001111101011101011010000010010111010011111011011001001110001111001101111011110010101010011010100110100010000001110111110000000101011001100001110001010110010110110010100010011000000001010011110110101100000110111100000100001111000100111100100101100111001101100001100011110110000100110111100010000001000101110001101111001101010011110 ;
  localparam Weights1 = 400'b1000001001011000001111101001101100001110001111001010000101111101010001111111000101111100001100010101000001100011101000110111111101010100011110011110101101101010110100000100000110101110001101100001000100001011111111100000010110110100110100100001000011110110000000101111000000001110011011100010000111100001101000101011101000000000000011110011011101011110110111100000110001101000011011011111010000010000 ;

  localparam SumL = $clog2(M+1);
  wire [SumL*C-1:0] sums;

  seqlego #(.N(N),.B(B),.M(M),.C(C),.Weights0(Weights0),.Weights1(Weights1)) layers (
    .clk(clk),
    .rst(rst),
    .data(data),
    .out(sums)
  );

  argmax #(.N(C),.I($clog2(C)),.K(SumL)) result (
     .inx(sums),
     .outimax(klass)
  );

endmodule
