`timescale 1us/1ns









module tbwinewhite_tnn1_tnnpar #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1000


)();
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
reg clk;
reg [FEAT_CNT*FEAT_BITS-1:0] features;
wire [$clog2(CLASS_CNT)-1:0] prediction;
wire [FEAT_CNT*FEAT_BITS-1:0] testcases [TEST_CNT-1:0];
parameter Nsperiod=5000;
localparam period=Nsperiod/500;


assign testcases[0] = 44'h24446225335;
assign testcases[1] = 44'h45825120334;
assign testcases[2] = 44'h54823222437;
assign testcases[3] = 44'h53737322325;
assign testcases[4] = 44'h53737322325;
assign testcases[5] = 44'h54823222437;
assign testcases[6] = 44'h45725222244;
assign testcases[7] = 44'h24446225335;
assign testcases[8] = 44'h45825120334;
assign testcases[9] = 44'h84724120427;
assign testcases[10] = 44'ha6412110437;
assign testcases[11] = 44'h46624111427;
assign testcases[12] = 44'h78722110426;
assign testcases[13] = 44'hb6c15320414;
assign testcases[14] = 44'h48446215657;
assign testcases[15] = 44'h96814110414;
assign testcases[16] = 44'h43823220064;
assign testcases[17] = 44'hc3912210594;
assign testcases[18] = 44'h96616110446;
assign testcases[19] = 44'h45735222144;
assign testcases[20] = 44'hc3912210594;
assign testcases[21] = 44'h82713111444;
assign testcases[22] = 44'h65b24220435;
assign testcases[23] = 44'h35526130196;
assign testcases[24] = 44'h55a25120434;
assign testcases[25] = 44'h65839322335;
assign testcases[26] = 44'h54b25220335;
assign testcases[27] = 44'h66a35222435;
assign testcases[28] = 44'h95715120536;
assign testcases[29] = 44'hb9614210345;
assign testcases[30] = 44'h56735122437;
assign testcases[31] = 44'h63b21020317;
assign testcases[32] = 44'h74723220336;
assign testcases[33] = 44'h35a24220314;
assign testcases[34] = 44'h63936124233;
assign testcases[35] = 44'hc4714130435;
assign testcases[36] = 44'h52825121254;
assign testcases[37] = 44'h81615220345;
assign testcases[38] = 44'h23745224435;
assign testcases[39] = 44'h23745224435;
assign testcases[40] = 44'h43626380424;
assign testcases[41] = 44'h42625381434;
assign testcases[42] = 44'h54636132345;
assign testcases[43] = 44'h46725220334;
assign testcases[44] = 44'h46825220324;
assign testcases[45] = 44'h56626220326;
assign testcases[46] = 44'h56827331364;
assign testcases[47] = 44'h56827331264;
assign testcases[48] = 44'h54636132345;
assign testcases[49] = 44'h55925231325;
assign testcases[50] = 44'ha4916230325;
assign testcases[51] = 44'h87914230334;
assign testcases[52] = 44'h74913120314;
assign testcases[53] = 44'h72914220324;
assign testcases[54] = 44'h33525270625;
assign testcases[55] = 44'h86617210335;
assign testcases[56] = 44'h45538223325;
assign testcases[57] = 44'h23835323323;
assign testcases[58] = 44'h63623121154;
assign testcases[59] = 44'h52924210326;
assign testcases[60] = 44'h24524241225;
assign testcases[61] = 44'h23835323323;
assign testcases[62] = 44'h62415110165;
assign testcases[63] = 44'h63623121154;
assign testcases[64] = 44'h64624210335;
assign testcases[65] = 44'h36724230044;
assign testcases[66] = 44'hc5714111234;
assign testcases[67] = 44'h54626420134;
assign testcases[68] = 44'h78923220324;
assign testcases[69] = 44'h42634122336;
assign testcases[70] = 44'h35639322434;
assign testcases[71] = 44'h47939321235;
assign testcases[72] = 44'h59e37231333;
assign testcases[73] = 44'h35322020427;
assign testcases[74] = 44'h78923220324;
assign testcases[75] = 44'h42634122336;
assign testcases[76] = 44'hc3813220325;
assign testcases[77] = 44'ha8912120345;
assign testcases[78] = 44'h36333132326;
assign testcases[79] = 44'h33824121374;
assign testcases[80] = 44'h7aa24220325;
assign testcases[81] = 44'h37746324325;
assign testcases[82] = 44'h54726331245;
assign testcases[83] = 44'h44937222325;
assign testcases[84] = 44'h24635323655;
assign testcases[85] = 44'h24635323665;
assign testcases[86] = 44'h24535323655;
assign testcases[87] = 44'h45737423335;
assign testcases[88] = 44'h24635323655;
assign testcases[89] = 44'h24635323665;
assign testcases[90] = 44'h24535323655;
assign testcases[91] = 44'h35639422434;
assign testcases[92] = 44'hc3815310335;
assign testcases[93] = 44'hc4815310325;
assign testcases[94] = 44'h94715310316;
assign testcases[95] = 44'h34539323335;
assign testcases[96] = 44'h25636124643;
assign testcases[97] = 44'h93313110337;
assign testcases[98] = 44'h51233012449;
assign testcases[99] = 44'h25636124643;
assign testcases[100] = 44'h34437323436;
assign testcases[101] = 44'h44a36322315;
assign testcases[102] = 44'h43936323223;
assign testcases[103] = 44'h34446224446;
assign testcases[104] = 44'h34437323436;
assign testcases[105] = 44'h32734223315;
assign testcases[106] = 44'h44a36322315;
assign testcases[107] = 44'h37646314325;
assign testcases[108] = 44'h37646314325;
assign testcases[109] = 44'h67827220345;
assign testcases[110] = 44'h23236332514;
assign testcases[111] = 44'h26549224435;
assign testcases[112] = 44'h35437423545;
assign testcases[113] = 44'h35735222354;
assign testcases[114] = 44'h35735222354;
assign testcases[115] = 44'h43d23030063;
assign testcases[116] = 44'h94915121243;
assign testcases[117] = 44'ha4713110415;
assign testcases[118] = 44'h35437423545;
assign testcases[119] = 44'h35537323545;
assign testcases[120] = 44'h65723121043;
assign testcases[121] = 44'h26435223336;
assign testcases[122] = 44'h42825222316;
assign testcases[123] = 44'h33825121325;
assign testcases[124] = 44'h53726240514;
assign testcases[125] = 44'h85815310324;
assign testcases[126] = 44'h64624212256;
assign testcases[127] = 44'h46b37312334;
assign testcases[128] = 44'h77826321534;
assign testcases[129] = 44'h77926221534;
assign testcases[130] = 44'h73a22012233;
assign testcases[131] = 44'h46b37312334;
assign testcases[132] = 44'h37739313454;
assign testcases[133] = 44'h35837214334;
assign testcases[134] = 44'h26737312235;
assign testcases[135] = 44'h46836214334;
assign testcases[136] = 44'h73624210427;
assign testcases[137] = 44'h24635322655;
assign testcases[138] = 44'h76613210325;
assign testcases[139] = 44'ha6723110437;
assign testcases[140] = 44'h64823120344;
assign testcases[141] = 44'h24635322655;
assign testcases[142] = 44'h76724210426;
assign testcases[143] = 44'h46723111427;
assign testcases[144] = 44'h86623110427;
assign testcases[145] = 44'h73414210434;
assign testcases[146] = 44'h53816320313;
assign testcases[147] = 44'h33a23121184;
assign testcases[148] = 44'ha7a13111344;
assign testcases[149] = 44'h43424121335;
assign testcases[150] = 44'h92625222426;
assign testcases[151] = 44'h54635322426;
assign testcases[152] = 44'h43424121335;
assign testcases[153] = 44'h64613220425;
assign testcases[154] = 44'h4c532122427;
assign testcases[155] = 44'h24237333436;
assign testcases[156] = 44'h24237333436;
assign testcases[157] = 44'hb4814210244;
assign testcases[158] = 44'hb2914210062;
assign testcases[159] = 44'hb2914210062;
assign testcases[160] = 44'hb4814210244;
assign testcases[161] = 44'h33436123524;
assign testcases[162] = 44'h73823121344;
assign testcases[163] = 44'h24237333436;
assign testcases[164] = 44'h45637323334;
assign testcases[165] = 44'h55636423325;
assign testcases[166] = 44'h47637222437;
assign testcases[167] = 44'hc4513110264;
assign testcases[168] = 44'h36535122336;
assign testcases[169] = 44'h51234012559;
assign testcases[170] = 44'hc6615230435;
assign testcases[171] = 44'h83613120426;
assign testcases[172] = 44'h93513010466;
assign testcases[173] = 44'h92914211424;
assign testcases[174] = 44'h68546224336;
assign testcases[175] = 44'h91625312425;
assign testcases[176] = 44'hc4512121545;
assign testcases[177] = 44'h43836323323;
assign testcases[178] = 44'h22624020193;
assign testcases[179] = 44'h39726221334;
assign testcases[180] = 44'h38726221344;
assign testcases[181] = 44'h34526320145;
assign testcases[182] = 44'h25346325435;
assign testcases[183] = 44'h47738323435;
assign testcases[184] = 44'h38438323535;
assign testcases[185] = 44'h38438423535;
assign testcases[186] = 44'h57636312434;
assign testcases[187] = 44'h85624211233;
assign testcases[188] = 44'hc7814111375;
assign testcases[189] = 44'h26537322334;
assign testcases[190] = 44'h26537322334;
assign testcases[191] = 44'h25346325435;
assign testcases[192] = 44'h93424122335;
assign testcases[193] = 44'h44924221314;
assign testcases[194] = 44'h34426491434;
assign testcases[195] = 44'h33426491434;
assign testcases[196] = 44'h33426491434;
assign testcases[197] = 44'h25638322235;
assign testcases[198] = 44'h25637323245;
assign testcases[199] = 44'h25638322235;
assign testcases[200] = 44'h35637324335;
assign testcases[201] = 44'h25637323245;
assign testcases[202] = 44'h45738323375;
assign testcases[203] = 44'ha6925213335;
assign testcases[204] = 44'h65824220333;
assign testcases[205] = 44'h24635223524;
assign testcases[206] = 44'h32734222315;
assign testcases[207] = 44'h5543412186a;
assign testcases[208] = 44'h6a923110385;
assign testcases[209] = 44'h4a726120354;
assign testcases[210] = 44'h62922112233;
assign testcases[211] = 44'h87914210425;
assign testcases[212] = 44'h32734222315;
assign testcases[213] = 44'h43a24221314;
assign testcases[214] = 44'h84814210234;
assign testcases[215] = 44'h43935322233;
assign testcases[216] = 44'h82526212336;
assign testcases[217] = 44'h43935322233;
assign testcases[218] = 44'h44946324233;
assign testcases[219] = 44'h82526212326;
assign testcases[220] = 44'h82526212336;
assign testcases[221] = 44'h36436232295;
assign testcases[222] = 44'h84814210234;
assign testcases[223] = 44'h33a25220324;
assign testcases[224] = 44'h66a25220274;
assign testcases[225] = 44'h23945224435;
assign testcases[226] = 44'h45b27220314;
assign testcases[227] = 44'h3673a422335;
assign testcases[228] = 44'h45b27220314;
assign testcases[229] = 44'h23945224435;
assign testcases[230] = 44'h24935132195;
assign testcases[231] = 44'h45937222437;
assign testcases[232] = 44'h45937312437;
assign testcases[233] = 44'h34537323425;
assign testcases[234] = 44'h34537323425;
assign testcases[235] = 44'h34537323425;
assign testcases[236] = 44'h34537323425;
assign testcases[237] = 44'h45838323375;
assign testcases[238] = 44'h84914210635;
assign testcases[239] = 44'h48b36114234;
assign testcases[240] = 44'h24747323245;
assign testcases[241] = 44'h65623112346;
assign testcases[242] = 44'h93613110425;
assign testcases[243] = 44'h47828321335;
assign testcases[244] = 44'h24635223555;
assign testcases[245] = 44'h9b929110324;
assign testcases[246] = 44'hc7615110325;
assign testcases[247] = 44'h73813110323;
assign testcases[248] = 44'h73812110323;
assign testcases[249] = 44'h54a34112154;
assign testcases[250] = 44'h59f37221323;
assign testcases[251] = 44'h55437234237;
assign testcases[252] = 44'h24635223555;
assign testcases[253] = 44'ha4c14011433;
assign testcases[254] = 44'h36726220433;
assign testcases[255] = 44'h47925210434;
assign testcases[256] = 44'h84823011344;
assign testcases[257] = 44'h84823011344;
assign testcases[258] = 44'ha5914110424;
assign testcases[259] = 44'h92812010443;
assign testcases[260] = 44'h64924221315;
assign testcases[261] = 44'h25345225435;
assign testcases[262] = 44'h62723112435;
assign testcases[263] = 44'h47538423435;
assign testcases[264] = 44'h75616110334;
assign testcases[265] = 44'h25345225435;
assign testcases[266] = 44'h35836222345;
assign testcases[267] = 44'h47925222182;
assign testcases[268] = 44'h47925222182;
assign testcases[269] = 44'h47925222182;
assign testcases[270] = 44'h35836222345;
assign testcases[271] = 44'h47925222182;
assign testcases[272] = 44'h33835223333;
assign testcases[273] = 44'h33824221384;
assign testcases[274] = 44'h47538322535;
assign testcases[275] = 44'h57636322424;
assign testcases[276] = 44'h57636322424;
assign testcases[277] = 44'h75212020436;
assign testcases[278] = 44'h75512120345;
assign testcases[279] = 44'hb9814111535;
assign testcases[280] = 44'hc3714111335;
assign testcases[281] = 44'hb7814211644;
assign testcases[282] = 44'h68527221465;
assign testcases[283] = 44'h35737324344;
assign testcases[284] = 44'h25647224245;
assign testcases[285] = 44'h25536322245;
assign testcases[286] = 44'h45737324334;
assign testcases[287] = 44'h35437323425;
assign testcases[288] = 44'h35437323425;
assign testcases[289] = 44'h35437323425;
assign testcases[290] = 44'h35437323425;
assign testcases[291] = 44'h64c25321313;
assign testcases[292] = 44'h34347335436;
assign testcases[293] = 44'h58a35122234;
assign testcases[294] = 44'h13736230488;
assign testcases[295] = 44'h46926220344;
assign testcases[296] = 44'h47536222757;
assign testcases[297] = 44'h87727421425;
assign testcases[298] = 44'h54735423416;
assign testcases[299] = 44'h64624120514;
assign testcases[300] = 44'h78813230054;
assign testcases[301] = 44'h63622120327;
assign testcases[302] = 44'h78813230054;
assign testcases[303] = 44'h84916220233;
assign testcases[304] = 44'h54726222255;
assign testcases[305] = 44'h54726222255;
assign testcases[306] = 44'h54726221255;
assign testcases[307] = 44'h54726221255;
assign testcases[308] = 44'h64725211344;
assign testcases[309] = 44'h64725211344;
assign testcases[310] = 44'h99a13110344;
assign testcases[311] = 44'hc5c16212172;
assign testcases[312] = 44'h54935221436;
assign testcases[313] = 44'h58826311243;
assign testcases[314] = 44'h57826311243;
assign testcases[315] = 44'h34524260635;
assign testcases[316] = 44'h73725211335;
assign testcases[317] = 44'h63725212334;
assign testcases[318] = 44'h94c25112533;
assign testcases[319] = 44'h57c22011214;
assign testcases[320] = 44'h67d22120203;
assign testcases[321] = 44'h63725212334;
assign testcases[322] = 44'h73725211335;
assign testcases[323] = 44'h63625212435;
assign testcases[324] = 44'h96427120557;
assign testcases[325] = 44'h6772b721336;
assign testcases[326] = 44'h57338214436;
assign testcases[327] = 44'h58725211244;
assign testcases[328] = 44'h45737324334;
assign testcases[329] = 44'h65723210425;
assign testcases[330] = 44'hc7913211344;
assign testcases[331] = 44'h73725211335;
assign testcases[332] = 44'ha3813110324;
assign testcases[333] = 44'h54635212334;
assign testcases[334] = 44'h73823111333;
assign testcases[335] = 44'ha3813110324;
assign testcases[336] = 44'h84914110324;
assign testcases[337] = 44'h34836323333;
assign testcases[338] = 44'h66b25120433;
assign testcases[339] = 44'h6ca25320324;
assign testcases[340] = 44'h36735122426;
assign testcases[341] = 44'h56724120336;
assign testcases[342] = 44'h35735222434;
assign testcases[343] = 44'h5a825221542;
assign testcases[344] = 44'h5a825321532;
assign testcases[345] = 44'h43825221315;
assign testcases[346] = 44'h85912110143;
assign testcases[347] = 44'h24745424424;
assign testcases[348] = 44'h55634223426;
assign testcases[349] = 44'h55635323416;
assign testcases[350] = 44'h9a815320314;
assign testcases[351] = 44'ha1525212445;
assign testcases[352] = 44'h45624130343;
assign testcases[353] = 44'ha1525212445;
assign testcases[354] = 44'h47829221453;
assign testcases[355] = 44'h33237333425;
assign testcases[356] = 44'h33237333425;
assign testcases[357] = 44'h4a626120344;
assign testcases[358] = 44'h6442512042a;
assign testcases[359] = 44'h77726211335;
assign testcases[360] = 44'h65836324334;
assign testcases[361] = 44'h24623120145;
assign testcases[362] = 44'h43a24221315;
assign testcases[363] = 44'h33237333425;
assign testcases[364] = 44'h94b23110415;
assign testcases[365] = 44'hb9a14211333;
assign testcases[366] = 44'h77b25240323;
assign testcases[367] = 44'h44625220245;
assign testcases[368] = 44'h78726220536;
assign testcases[369] = 44'h91722123355;
assign testcases[370] = 44'h44625220245;
assign testcases[371] = 44'h78726220536;
assign testcases[372] = 44'h569271202d4;
assign testcases[373] = 44'h35625220335;
assign testcases[374] = 44'hc3b13110242;
assign testcases[375] = 44'hc3b13110242;
assign testcases[376] = 44'h65914110344;
assign testcases[377] = 44'h54623120425;
assign testcases[378] = 44'h58725120543;
assign testcases[379] = 44'h65914110344;
assign testcases[380] = 44'h54623120425;
assign testcases[381] = 44'h36636323335;
assign testcases[382] = 44'h36635122346;
assign testcases[383] = 44'h35625220335;
assign testcases[384] = 44'h93a14111443;
assign testcases[385] = 44'hc3b13110242;
assign testcases[386] = 44'h73b14110512;
assign testcases[387] = 44'h58629411354;
assign testcases[388] = 44'h44a25221324;
assign testcases[389] = 44'h37736314435;
assign testcases[390] = 44'h37736314435;
assign testcases[391] = 44'h74612110344;
assign testcases[392] = 44'h65934112174;
assign testcases[393] = 44'hb6512110435;
assign testcases[394] = 44'h24736323555;
assign testcases[395] = 44'h54726510135;
assign testcases[396] = 44'h93513210437;
assign testcases[397] = 44'h95b14210424;
assign testcases[398] = 44'h44946324333;
assign testcases[399] = 44'ha4813211424;
assign testcases[400] = 44'h95b14210424;
assign testcases[401] = 44'h24736323555;
assign testcases[402] = 44'h36724130144;
assign testcases[403] = 44'h26549324335;
assign testcases[404] = 44'hc8816211325;
assign testcases[405] = 44'h54726510135;
assign testcases[406] = 44'hc3a13211333;
assign testcases[407] = 44'h45724120265;
assign testcases[408] = 44'h66824120414;
assign testcases[409] = 44'h93513210437;
assign testcases[410] = 44'h35445215435;
assign testcases[411] = 44'h4b835213335;
assign testcases[412] = 44'h65613210425;
assign testcases[413] = 44'h65613210425;
assign testcases[414] = 44'h35445215435;
assign testcases[415] = 44'h4b835213335;
assign testcases[416] = 44'h52723120326;
assign testcases[417] = 44'h35637322235;
assign testcases[418] = 44'h52723120326;
assign testcases[419] = 44'h66925220346;
assign testcases[420] = 44'hc3615211325;
assign testcases[421] = 44'h66838222325;
assign testcases[422] = 44'h66838222325;
assign testcases[423] = 44'h66838222325;
assign testcases[424] = 44'h66936322425;
assign testcases[425] = 44'h66838222325;
assign testcases[426] = 44'h66838222325;
assign testcases[427] = 44'h44537323535;
assign testcases[428] = 44'h34523120326;
assign testcases[429] = 44'h35637323545;
assign testcases[430] = 44'h44537323535;
assign testcases[431] = 44'h53723120144;
assign testcases[432] = 44'h57728420316;
assign testcases[433] = 44'h37525150175;
assign testcases[434] = 44'hb5924212325;
assign testcases[435] = 44'hb5a23111425;
assign testcases[436] = 44'h57828120334;
assign testcases[437] = 44'hb8917310314;
assign testcases[438] = 44'h57728420316;
assign testcases[439] = 44'h36824120044;
assign testcases[440] = 44'h97813110424;
assign testcases[441] = 44'h69825111254;
assign testcases[442] = 44'hd8a14310333;
assign testcases[443] = 44'h36839323474;
assign testcases[444] = 44'h82735215335;
assign testcases[445] = 44'h93822113345;
assign testcases[446] = 44'hb4c15220333;
assign testcases[447] = 44'h56a34123254;
assign testcases[448] = 44'h56a34123254;
assign testcases[449] = 44'h66b24220334;
assign testcases[450] = 44'h36536132285;
assign testcases[451] = 44'h54824210224;
assign testcases[452] = 44'h75b26121163;
assign testcases[453] = 44'h65a24220333;
assign testcases[454] = 44'h66b24220334;
assign testcases[455] = 44'h56a34123254;
assign testcases[456] = 44'hd3813110324;
assign testcases[457] = 44'h46334122325;
assign testcases[458] = 44'h59828220353;
assign testcases[459] = 44'h15939522354;
assign testcases[460] = 44'h46334122325;
assign testcases[461] = 44'h34736224335;
assign testcases[462] = 44'h43936323233;
assign testcases[463] = 44'h43722120245;
assign testcases[464] = 44'h25636423655;
assign testcases[465] = 44'h24334232624;
assign testcases[466] = 44'h44735312315;
assign testcases[467] = 44'h43722120245;
assign testcases[468] = 44'h25636423655;
assign testcases[469] = 44'h46546324535;
assign testcases[470] = 44'h39436113757;
assign testcases[471] = 44'h5a627211354;
assign testcases[472] = 44'hc4813110334;
assign testcases[473] = 44'h45925211315;
assign testcases[474] = 44'h43823211213;
assign testcases[475] = 44'h47538313535;
assign testcases[476] = 44'hb3414210336;
assign testcases[477] = 44'h66624210325;
assign testcases[478] = 44'h37426130175;
assign testcases[479] = 44'h66926420324;
assign testcases[480] = 44'h37736222364;
assign testcases[481] = 44'h75914220443;
assign testcases[482] = 44'h44935223233;
assign testcases[483] = 44'h37736222364;
assign testcases[484] = 44'h478374f1354;
assign testcases[485] = 44'h46b24210424;
assign testcases[486] = 44'h45b24210413;
assign testcases[487] = 44'h74613210344;
assign testcases[488] = 44'h69926320336;
assign testcases[489] = 44'h24636322336;
assign testcases[490] = 44'hb4512010335;
assign testcases[491] = 44'hc3812110425;
assign testcases[492] = 44'h54736212326;
assign testcases[493] = 44'h98716110324;
assign testcases[494] = 44'h77923111425;
assign testcases[495] = 44'hc5916112163;
assign testcases[496] = 44'h25537423655;
assign testcases[497] = 44'hc6815210325;
assign testcases[498] = 44'h58826110343;
assign testcases[499] = 44'h25537423655;
assign testcases[500] = 44'h45547324535;
assign testcases[501] = 44'h45636313625;
assign testcases[502] = 44'h57727010334;
assign testcases[503] = 44'h57727010334;
assign testcases[504] = 44'h26535223326;
assign testcases[505] = 44'h26535223326;
assign testcases[506] = 44'h26425041375;
assign testcases[507] = 44'h56d26220333;
assign testcases[508] = 44'ha4a15311383;
assign testcases[509] = 44'h56d26220333;
assign testcases[510] = 44'h54725320134;
assign testcases[511] = 44'hb4616020346;
assign testcases[512] = 44'h87625211335;
assign testcases[513] = 44'h82712110346;
assign testcases[514] = 44'h63724212336;
assign testcases[515] = 44'h65926120344;
assign testcases[516] = 44'h34525320425;
assign testcases[517] = 44'h67425320416;
assign testcases[518] = 44'h78a13120313;
assign testcases[519] = 44'ha3721023345;
assign testcases[520] = 44'h5a525010326;
assign testcases[521] = 44'h5a525010326;
assign testcases[522] = 44'h93513110435;
assign testcases[523] = 44'h83513110343;
assign testcases[524] = 44'h92912010443;
assign testcases[525] = 44'h34525151443;
assign testcases[526] = 44'hc6511011445;
assign testcases[527] = 44'hc4914210234;
assign testcases[528] = 44'hb2a14110042;
assign testcases[529] = 44'h84c24111523;
assign testcases[530] = 44'h4ba23221304;
assign testcases[531] = 44'h33525381524;
assign testcases[532] = 44'h35436333336;
assign testcases[533] = 44'h35436333336;
assign testcases[534] = 44'h35436333336;
assign testcases[535] = 44'h35546324546;
assign testcases[536] = 44'h35546324546;
assign testcases[537] = 44'h35436333336;
assign testcases[538] = 44'h66922120334;
assign testcases[539] = 44'h48937221235;
assign testcases[540] = 44'h96b36012344;
assign testcases[541] = 44'h24637422665;
assign testcases[542] = 44'h59926120343;
assign testcases[543] = 44'h57725212434;
assign testcases[544] = 44'h35736323235;
assign testcases[545] = 44'h57b25210214;
assign testcases[546] = 44'h48b36212234;
assign testcases[547] = 44'ha5823020426;
assign testcases[548] = 44'h65b24220324;
assign testcases[549] = 44'h24637422665;
assign testcases[550] = 44'h46536223535;
assign testcases[551] = 44'h93313210338;
assign testcases[552] = 44'hb3414210336;
assign testcases[553] = 44'h46536223535;
assign testcases[554] = 44'hb3414210336;
assign testcases[555] = 44'h93313210338;
assign testcases[556] = 44'h48436123747;
assign testcases[557] = 44'h65925120254;
assign testcases[558] = 44'h43836323223;
assign testcases[559] = 44'hba415321445;
assign testcases[560] = 44'h5a635222424;
assign testcases[561] = 44'h55824220153;
assign testcases[562] = 44'h38536232346;
assign testcases[563] = 44'h6a525120236;
assign testcases[564] = 44'h34726231375;
assign testcases[565] = 44'h55633122426;
assign testcases[566] = 44'h93621023345;
assign testcases[567] = 44'h57525320533;
assign testcases[568] = 44'h57525320534;
assign testcases[569] = 44'h49726211334;
assign testcases[570] = 44'h24537423656;
assign testcases[571] = 44'h94914111334;
assign testcases[572] = 44'h26546224544;
assign testcases[573] = 44'hc3615311325;
assign testcases[574] = 44'ha4715210326;
assign testcases[575] = 44'h65627320327;
assign testcases[576] = 44'h65627320327;
assign testcases[577] = 44'hc3615311325;
assign testcases[578] = 44'h94914111334;
assign testcases[579] = 44'hb3a15211353;
assign testcases[580] = 44'h24537423656;
assign testcases[581] = 44'h43924121223;
assign testcases[582] = 44'h52626221235;
assign testcases[583] = 44'h43233122236;
assign testcases[584] = 44'h55a25220334;
assign testcases[585] = 44'h43233122236;
assign testcases[586] = 44'h25635222336;
assign testcases[587] = 44'h75b25210244;
assign testcases[588] = 44'h75a24210335;
assign testcases[589] = 44'h47725111325;
assign testcases[590] = 44'h34335023545;
assign testcases[591] = 44'h75924310425;
assign testcases[592] = 44'h46735122355;
assign testcases[593] = 44'h71415010164;
assign testcases[594] = 44'h71415010164;
assign testcases[595] = 44'h65b25020434;
assign testcases[596] = 44'h46735122355;
assign testcases[597] = 44'h74724111435;
assign testcases[598] = 44'h65924213333;
assign testcases[599] = 44'h99512110425;
assign testcases[600] = 44'h46626280334;
assign testcases[601] = 44'h73214220435;
assign testcases[602] = 44'h71415010164;
assign testcases[603] = 44'h71415010164;
assign testcases[604] = 44'h57425220534;
assign testcases[605] = 44'h57425220534;
assign testcases[606] = 44'h43a36222335;
assign testcases[607] = 44'h43a36222335;
assign testcases[608] = 44'h45946324234;
assign testcases[609] = 44'h79b33121356;
assign testcases[610] = 44'hb8814211344;
assign testcases[611] = 44'h83523011436;
assign testcases[612] = 44'h23435223726;
assign testcases[613] = 44'h23435223726;
assign testcases[614] = 44'h23435223726;
assign testcases[615] = 44'h23435223726;
assign testcases[616] = 44'ha8713110346;
assign testcases[617] = 44'h75727320336;
assign testcases[618] = 44'h75727320336;
assign testcases[619] = 44'h45625220326;
assign testcases[620] = 44'h37748344464;
assign testcases[621] = 44'h35236342434;
assign testcases[622] = 44'h67925121142;
assign testcases[623] = 44'h95712020335;
assign testcases[624] = 44'h36824130143;
assign testcases[625] = 44'h84924313334;
assign testcases[626] = 44'h34936142186;
assign testcases[627] = 44'h47738221245;
assign testcases[628] = 44'h47738221245;
assign testcases[629] = 44'h67713110343;
assign testcases[630] = 44'h24745224425;
assign testcases[631] = 44'h24745224425;
assign testcases[632] = 44'h78825111335;
assign testcases[633] = 44'h44937223233;
assign testcases[634] = 44'h75a25211314;
assign testcases[635] = 44'h75b25211213;
assign testcases[636] = 44'h74a25211314;
assign testcases[637] = 44'h37635123236;
assign testcases[638] = 44'h69827321143;
assign testcases[639] = 44'h69827321143;
assign testcases[640] = 44'h85914220323;
assign testcases[641] = 44'h34837223234;
assign testcases[642] = 44'h65936423324;
assign testcases[643] = 44'h44936223334;
assign testcases[644] = 44'h44936223334;
assign testcases[645] = 44'h34836222234;
assign testcases[646] = 44'h47525020744;
assign testcases[647] = 44'h33635323306;
assign testcases[648] = 44'h59627221143;
assign testcases[649] = 44'h36547233335;
assign testcases[650] = 44'h36547233335;
assign testcases[651] = 44'h36547233335;
assign testcases[652] = 44'h36547233335;
assign testcases[653] = 44'h44935223333;
assign testcases[654] = 44'h9a915420424;
assign testcases[655] = 44'hb4624211336;
assign testcases[656] = 44'h93523111338;
assign testcases[657] = 44'h64825121245;
assign testcases[658] = 44'h93817221234;
assign testcases[659] = 44'h55628710235;
assign testcases[660] = 44'h43623120335;
assign testcases[661] = 44'hb5925313335;
assign testcases[662] = 44'h35a37142185;
assign testcases[663] = 44'h43623120335;
assign testcases[664] = 44'h46936322415;
assign testcases[665] = 44'h45824120236;
assign testcases[666] = 44'hc9917210425;
assign testcases[667] = 44'h46936322415;
assign testcases[668] = 44'h54926220214;
assign testcases[669] = 44'h37737323534;
assign testcases[670] = 44'h36637222356;
assign testcases[671] = 44'h97813110334;
assign testcases[672] = 44'hc5a25213345;
assign testcases[673] = 44'h78924110344;
assign testcases[674] = 44'h47537322544;
assign testcases[675] = 44'h33737222234;
assign testcases[676] = 44'h34738323233;
assign testcases[677] = 44'ha4a13111443;
assign testcases[678] = 44'ha4a13111443;
assign testcases[679] = 44'ha4a13111443;
assign testcases[680] = 44'h53726320134;
assign testcases[681] = 44'h45526120745;
assign testcases[682] = 44'h44836223233;
assign testcases[683] = 44'h456263b1334;
assign testcases[684] = 44'h84526320367;
assign testcases[685] = 44'h34837323344;
assign testcases[686] = 44'h76824121325;
assign testcases[687] = 44'h385371d3395;
assign testcases[688] = 44'h35638322335;
assign testcases[689] = 44'h77824210414;
assign testcases[690] = 44'h57925120325;
assign testcases[691] = 44'h57727211244;
assign testcases[692] = 44'h57727211243;
assign testcases[693] = 44'h58727211153;
assign testcases[694] = 44'h48648324636;
assign testcases[695] = 44'h44737323344;
assign testcases[696] = 44'h87713110324;
assign testcases[697] = 44'h47537313546;
assign testcases[698] = 44'h47537313546;
assign testcases[699] = 44'h47537323546;
assign testcases[700] = 44'h48537223757;
assign testcases[701] = 44'hfaa15110243;
assign testcases[702] = 44'h54723120254;
assign testcases[703] = 44'h64614210344;
assign testcases[704] = 44'hc5a14111333;
assign testcases[705] = 44'h72221111437;
assign testcases[706] = 44'h57628321244;
assign testcases[707] = 44'h87626321425;
assign testcases[708] = 44'h55644223426;
assign testcases[709] = 44'h34623120264;
assign testcases[710] = 44'h44936323234;
assign testcases[711] = 44'hb5614210437;
assign testcases[712] = 44'hb5614210437;
assign testcases[713] = 44'h54928312444;
assign testcases[714] = 44'h75a27211353;
assign testcases[715] = 44'h69b25210324;
assign testcases[716] = 44'h37538122356;
assign testcases[717] = 44'h35345224435;
assign testcases[718] = 44'h69b25210324;
assign testcases[719] = 44'h65b24220536;
assign testcases[720] = 44'h24436322434;
assign testcases[721] = 44'h66b26120433;
assign testcases[722] = 44'ha5914110345;
assign testcases[723] = 44'hb4813210344;
assign testcases[724] = 44'h73614110436;
assign testcases[725] = 44'h64625220254;
assign testcases[726] = 44'ha8914211334;
assign testcases[727] = 44'h47433122325;
assign testcases[728] = 44'h65925221314;
assign testcases[729] = 44'h47627180343;
assign testcases[730] = 44'h66935123324;
assign testcases[731] = 44'h45839422534;
assign testcases[732] = 44'h82421111438;
assign testcases[733] = 44'h35436223334;
assign testcases[734] = 44'h37837112255;
assign testcases[735] = 44'h45624111334;
assign testcases[736] = 44'h35436223334;
assign testcases[737] = 44'h37837112255;
assign testcases[738] = 44'h73725211325;
assign testcases[739] = 44'h45624111334;
assign testcases[740] = 44'hc3910011455;
assign testcases[741] = 44'h86a12110323;
assign testcases[742] = 44'h67825110425;
assign testcases[743] = 44'h44935213233;
assign testcases[744] = 44'h54736122356;
assign testcases[745] = 44'hb6814210f26;
assign testcases[746] = 44'h66739212325;
assign testcases[747] = 44'h92526312435;
assign testcases[748] = 44'h56836222425;
assign testcases[749] = 44'h92526312435;
assign testcases[750] = 44'h92526312435;
assign testcases[751] = 44'h66636412525;
assign testcases[752] = 44'h45646513424;
assign testcases[753] = 44'h66739212325;
assign testcases[754] = 44'h35525150543;
assign testcases[755] = 44'hb5814210435;
assign testcases[756] = 44'h44a36223333;
assign testcases[757] = 44'h3ca46424425;
assign testcases[758] = 44'h5e825320415;
assign testcases[759] = 44'h5e825320415;
assign testcases[760] = 44'h56836222425;
assign testcases[761] = 44'h56836222425;
assign testcases[762] = 44'h26449325535;
assign testcases[763] = 44'h67944214062;
assign testcases[764] = 44'h49726221334;
assign testcases[765] = 44'h84325220435;
assign testcases[766] = 44'h34549433674;
assign testcases[767] = 44'h77711010325;
assign testcases[768] = 44'h33a34222304;
assign testcases[769] = 44'h33a34222304;
assign testcases[770] = 44'h54a24221315;
assign testcases[771] = 44'h33625360514;
assign testcases[772] = 44'h33625360624;
assign testcases[773] = 44'h44a46314334;
assign testcases[774] = 44'h64734112438;
assign testcases[775] = 44'hb7814250524;
assign testcases[776] = 44'h86423110417;
assign testcases[777] = 44'h36647323225;
assign testcases[778] = 44'h4b946324425;
assign testcases[779] = 44'h2a845223417;
assign testcases[780] = 44'h83912020053;
assign testcases[781] = 44'h37538222236;
assign testcases[782] = 44'h4b946324425;
assign testcases[783] = 44'h2a845223417;
assign testcases[784] = 44'h36647323225;
assign testcases[785] = 44'h31834212336;
assign testcases[786] = 44'h31834213346;
assign testcases[787] = 44'h31834213346;
assign testcases[788] = 44'h54b24112243;
assign testcases[789] = 44'h31834212336;
assign testcases[790] = 44'h31834213346;
assign testcases[791] = 44'h79a23110333;
assign testcases[792] = 44'h56625221164;
assign testcases[793] = 44'h79a23110333;
assign testcases[794] = 44'h36526220346;
assign testcases[795] = 44'h34535222345;
assign testcases[796] = 44'h37438222256;
assign testcases[797] = 44'h4a835323335;
assign testcases[798] = 44'h43a24221222;
assign testcases[799] = 44'h87912110323;
assign testcases[800] = 44'h24536213636;
assign testcases[801] = 44'h35738322533;
assign testcases[802] = 44'h36538323355;
assign testcases[803] = 44'h54a36213324;
assign testcases[804] = 44'h54724111345;
assign testcases[805] = 44'h24536213636;
assign testcases[806] = 44'h44737323344;
assign testcases[807] = 44'h44637323334;
assign testcases[808] = 44'h33639423253;
assign testcases[809] = 44'h44737323334;
assign testcases[810] = 44'h35738322533;
assign testcases[811] = 44'h36724130053;
assign testcases[812] = 44'h35a26020344;
assign testcases[813] = 44'h44a46224334;
assign testcases[814] = 44'h67538234246;
assign testcases[815] = 44'h34424111234;
assign testcases[816] = 44'ha6623011427;
assign testcases[817] = 44'h35735112284;
assign testcases[818] = 44'h34424111234;
assign testcases[819] = 44'h35735112284;
assign testcases[820] = 44'hb7a13110344;
assign testcases[821] = 44'h37338132295;
assign testcases[822] = 44'h44824221225;
assign testcases[823] = 44'h44924221224;
assign testcases[824] = 44'ha6623011427;
assign testcases[825] = 44'h56836222425;
assign testcases[826] = 44'h67935122435;
assign testcases[827] = 44'hc5815110336;
assign testcases[828] = 44'h74633122315;
assign testcases[829] = 44'h84623120315;
assign testcases[830] = 44'h69f34220325;
assign testcases[831] = 44'h97526211416;
assign testcases[832] = 44'hc6914221335;
assign testcases[833] = 44'hb4713110335;
assign testcases[834] = 44'h69f34220325;
assign testcases[835] = 44'hc4614211356;
assign testcases[836] = 44'ha3816210335;
assign testcases[837] = 44'ha3816210335;
assign testcases[838] = 44'ha3816210335;
assign testcases[839] = 44'ha3624111346;
assign testcases[840] = 44'ha3624111346;
assign testcases[841] = 44'h25646223328;
assign testcases[842] = 44'h25646223328;
assign testcases[843] = 44'h76723210325;
assign testcases[844] = 44'h85814210325;
assign testcases[845] = 44'h85814210325;
assign testcases[846] = 44'h33435314424;
assign testcases[847] = 44'h73522110348;
assign testcases[848] = 44'h25646223328;
assign testcases[849] = 44'h95914210223;
assign testcases[850] = 44'h76723210325;
assign testcases[851] = 44'h46646323557;
assign testcases[852] = 44'h4e824210325;
assign testcases[853] = 44'h25535213646;
assign testcases[854] = 44'h4e824210325;
assign testcases[855] = 44'h6ab24210326;
assign testcases[856] = 44'h46646323557;
assign testcases[857] = 44'h46646323557;
assign testcases[858] = 44'h56735312424;
assign testcases[859] = 44'h45726381334;
assign testcases[860] = 44'h68723210337;
assign testcases[861] = 44'h3a846323435;
assign testcases[862] = 44'h57926211042;
assign testcases[863] = 44'hb5814110334;
assign testcases[864] = 44'h57926211042;
assign testcases[865] = 44'hc1604110334;
assign testcases[866] = 44'h4e824210325;
assign testcases[867] = 44'h1a845223426;
assign testcases[868] = 44'h3b846313435;
assign testcases[869] = 44'h59723210335;
assign testcases[870] = 44'h45536132663;
assign testcases[871] = 44'h25535213646;
assign testcases[872] = 44'h72514111234;
assign testcases[873] = 44'h4122101051a;
assign testcases[874] = 44'h53922010316;
assign testcases[875] = 44'h57725110325;
assign testcases[876] = 44'hc3814301345;
assign testcases[877] = 44'h63724250333;
assign testcases[878] = 44'h23724260514;
assign testcases[879] = 44'haba14110315;
assign testcases[880] = 44'h57725110325;
assign testcases[881] = 44'h55734010448;
assign testcases[882] = 44'h96624111436;
assign testcases[883] = 44'h96624111436;
assign testcases[884] = 44'h56938213325;
assign testcases[885] = 44'hb8a14110344;
assign testcases[886] = 44'h95716210335;
assign testcases[887] = 44'h89913220334;
assign testcases[888] = 44'h95716210335;
assign testcases[889] = 44'h89913220334;
assign testcases[890] = 44'h58826221042;
assign testcases[891] = 44'h83a14210233;
assign testcases[892] = 44'h45d24210333;
assign testcases[893] = 44'hb3614210345;
assign testcases[894] = 44'h83a14210233;
assign testcases[895] = 44'h66712120423;
assign testcases[896] = 44'h66729322325;
assign testcases[897] = 44'h64523120335;
assign testcases[898] = 44'h75512110334;
assign testcases[899] = 44'h66729322325;
assign testcases[900] = 44'h86925222424;
assign testcases[901] = 44'h43834123336;
assign testcases[902] = 44'h23538323334;
assign testcases[903] = 44'h43727322343;
assign testcases[904] = 44'h25426320325;
assign testcases[905] = 44'h88523020427;
assign testcases[906] = 44'h67522020437;
assign testcases[907] = 44'hb4814210435;
assign testcases[908] = 44'h55936122426;
assign testcases[909] = 44'h26548223336;
assign testcases[910] = 44'h58625111244;
assign testcases[911] = 44'h58625121244;
assign testcases[912] = 44'h58625121244;
assign testcases[913] = 44'h32921110033;
assign testcases[914] = 44'h43823120346;
assign testcases[915] = 44'h32921110033;
assign testcases[916] = 44'h66925221416;
assign testcases[917] = 44'h82314110336;
assign testcases[918] = 44'ha3514110335;
assign testcases[919] = 44'h62324110427;
assign testcases[920] = 44'h44c35321305;
assign testcases[921] = 44'h24635312646;
assign testcases[922] = 44'h24635312646;
assign testcases[923] = 44'h54738423334;
assign testcases[924] = 44'h75b25320436;
assign testcases[925] = 44'h54823121234;
assign testcases[926] = 44'h33923121182;
assign testcases[927] = 44'h45426321334;
assign testcases[928] = 44'h55d36323334;
assign testcases[929] = 44'h35634224644;
assign testcases[930] = 44'ha3623101516;
assign testcases[931] = 44'h23538313434;
assign testcases[932] = 44'h54738423334;
assign testcases[933] = 44'h44827312333;
assign testcases[934] = 44'h23538313434;
assign testcases[935] = 44'h23628321434;
assign testcases[936] = 44'h94522020354;
assign testcases[937] = 44'h35634224644;
assign testcases[938] = 44'h56939322344;
assign testcases[939] = 44'h45537224336;
assign testcases[940] = 44'h47627212344;
assign testcases[941] = 44'h46838313434;
assign testcases[942] = 44'h54c23110252;
assign testcases[943] = 44'hb3615211365;
assign testcases[944] = 44'h24835122324;
assign testcases[945] = 44'h64c24121314;
assign testcases[946] = 44'h44347324a47;
assign testcases[947] = 44'h53325110317;
assign testcases[948] = 44'h469320212a5;
assign testcases[949] = 44'h94723011435;
assign testcases[950] = 44'h43525120346;
assign testcases[951] = 44'h55535112326;
assign testcases[952] = 44'h56723110314;
assign testcases[953] = 44'h53424220427;
assign testcases[954] = 44'h55535112326;
assign testcases[955] = 44'h43525120346;
assign testcases[956] = 44'h43525120346;
assign testcases[957] = 44'h66a23120324;
assign testcases[958] = 44'h66a23110324;
assign testcases[959] = 44'h34536224335;
assign testcases[960] = 44'h34536224335;
assign testcases[961] = 44'hb7623211356;
assign testcases[962] = 44'h34536224335;
assign testcases[963] = 44'h95924111224;
assign testcases[964] = 44'h44835213233;
assign testcases[965] = 44'h93623111427;
assign testcases[966] = 44'h43627220344;
assign testcases[967] = 44'h34845214325;
assign testcases[968] = 44'ha9913110304;
assign testcases[969] = 44'h95912100153;
assign testcases[970] = 44'hb3a13100052;
assign testcases[971] = 44'hc5914110233;
assign testcases[972] = 44'h34845214325;
assign testcases[973] = 44'ha9913110304;
assign testcases[974] = 44'had924120415;
assign testcases[975] = 44'h35634121236;
assign testcases[976] = 44'h64b25321314;
assign testcases[977] = 44'h25837322314;
assign testcases[978] = 44'h77a25211336;
assign testcases[979] = 44'h55622070723;
assign testcases[980] = 44'h54622070723;
assign testcases[981] = 44'h77a25211336;
assign testcases[982] = 44'hc4b12110252;
assign testcases[983] = 44'ha4a13111343;
assign testcases[984] = 44'h76a25320325;
assign testcases[985] = 44'h66a24220253;
assign testcases[986] = 44'h65626221336;
assign testcases[987] = 44'h64626221336;
assign testcases[988] = 44'h76a25320325;
assign testcases[989] = 44'ha3524012436;
assign testcases[990] = 44'h63325211417;
assign testcases[991] = 44'h67622020437;
assign testcases[992] = 44'h53738424334;
assign testcases[993] = 44'h55a22020235;
assign testcases[994] = 44'h46837110327;
assign testcases[995] = 44'h64525120336;
assign testcases[996] = 44'h68821020333;
assign testcases[997] = 44'h45935232334;
assign testcases[998] = 44'h35546224336;
assign testcases[999] = 44'h56526320626;



winewhite_tnn1_tnnpar dut (.features(features),.prediction(prediction));

integer i,j;
initial begin
    features = testcases[0];
    for(i=0;i<TEST_CNT;i=i+1) begin
        features = testcases[i];
        #period
        for(j=0;j<CLASS_CNT;j=j+1) begin
            $write("%d ,",dut.scores[j]);
        end
        $display("");
    end
end

endmodule
