
















module pendigits_tnn1_tnnpaarter #(

parameter FEAT_CNT = 16,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 10,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 7584'h0005008a0001001400890001001f00880001001c00870001005f00850001000d00840001001d00830001000b008200010022007f0001002b007e0001002b007d00010030007c00010079007b0001000e007a0001004200780001006a00770001000400760001002400740001000000730001004c007200010025006e00010048006d00010046006c0001002a006b0001000100690001005b00680001001c00660001004a006500010055006400010039006200010059005d00010042005a0001003100560001001700470001000700370001005700710000005400700000003f006f00000035006700000032006300000032006100000040006000000033005e00000036005c0000003e00580000002900530000001900520000002d005100000035005000000020004f0000003b004e00000036004d0000003f004b0000002c00490000001e00450000003d00440000003b00430000000c00430000003c00410000000900410000002800400000002b003e00000020003d00000027003c00000005003a0000001700390000001d00340000001700340000002c003300000015003100000014003000000027002f0000000d002f00000023002e00000023002d00000005002d0000000e002c0000002000270000000c00260000001600240000000500220000001900210000001300210000001a002000000008002000000015001f00000018001d0000000a001c00000019001b00000012001b0000000c001b00000004001600000003001500000009001300000000001000000002000f00000001000900000001000200000001000d00000004000c00000007000b00000004000a00000007000800000002000400000001000300000007003700000021002e0001001e002600010018001a0001000e001500010011001b00000011001300010005000600010024003800000003002a0000001200290000001c002800000008002300000009002200000010001c0000000a001700000008001600000004001500000003001300000009001a0001000200040001000b00190000001a001e0001001d00250001000d001f00010006001600010007000c00010017001900000001001400000004000f00000016001b0001000a000e00010001001400010002000c00010012001700010004001600010003001300010009000f0000000000060001000b001000000006001500010008001800000010001100000013001400000004000a00010010001100010002000500000008001200010003000900010001000700010000000c0000000b000e0000000d000f0000 ;
localparam YMAP = 1280'h0001008f000000a5000000a80001009500000096000100810000009e0001009f000100ab000100a600010097000000a70001009b000000ac000000800000009a000000ad00010093000000a10000003a0000009800000092000100a9000000aa0001008b0001008e0001008c000100900000009900010094000100750001009d000000860001008d000000a3000000a2000000910001009c000100a0000100a4;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 400'b0000000111000000011000100000000001001000000001010101101010000101011000000000000000000000000110101010000001010000000101000000000000000011000111010000110011100010100000000100010101000010010000001000001010001010101110000010000010001100000010000000000000000000110010001001001001010110100000000000001010000000110110010001010100000011000000001000001011010001000000000000000000001000000010000000010010001010 ;
localparam WNNZ = 400'b0010000111000010111010111001000011111000101011010111111110100111111010010101000000010000101110111010000001010000110111010010010100001011111111111101110111100010100010001100010101000010110101101000011110001011111111001111101011101100001011000000000011110000111010001101011101111111100000000101001010011000111110011111111100001011000101001100111011010111111000111000000100101001110011100101110110111110;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
wire [SUM_BITS-1:0] scorarr [CLASS_CNT-1:0];
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;

generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam adsub = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(adsub)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] <= 0;
end
endgenerate

function [7:0] zerocnt(input integer k);
    integer i,j;
    reg [HIDDEN_CNT-1:0] neur1;
    begin
        i = 0;
        neur1 = WNNZ[k*HIDDEN_CNT+:HIDDEN_CNT];
        for(j=0;j<HIDDEN_CNT;j=j+1)
            i = i + !(neur1[j]);
        zerocnt = i;
    end
endfunction

function [7:0] minzc(input integer k);
    integer i,j,h;
    begin
        i = HIDDEN_CNT;
        for(j=0;j<CLASS_CNT;j=j+1) begin
            h = zerocnt(j);
            if(h<i)
                i = h;
        end
        minzc = i;
    end
endfunction

localparam MINZC = minzc(0);

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    localparam Wuse = WNNZ[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wuse[j]) begin
            if(Wneur[j])
                tmpscore = tmpscore + hidden[j];
            else 
                tmpscore = tmpscore + hidden_n[j];
        end
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = 2*tmpscore + zerocnt(i) - MINZC;
    /* assign scorarr[i] = 2*tmpscore + zerocnt(i) - MINZC; */
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
