
















module cardio_tnn1_tnnpaarter #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 8832'h004500a40001005d00a30001000c00a20001009c00a10001003800a00001001b009f00010011009e0001002c009d00010095009b00010072009a0001007500990001008a00980001005a00970001000600960001008f00940001006200930001005c00920001007b009100010061009000010021008e00010078008d00010080008c0001002600890001006500880001001d00870001000700850001007c00830001003e008100010006007f00010017007e0001003d007a0001006a00790001003900770001005e00740001006d006f00010006006c0001004800640001001e002300010063008b0000005f00860000005600820000006000760000003300730000003400710000003f007000000043006e0000003b006b0000002600690000002c00680000003900670000004e006600000046005b0000002500590000003e00580000003000570000002d00550000001600540000001100530000002e00520000003200510000003d005000000026004f0000001c004d0000001e004c0000002b004b00000005004a0000003700490000002b004700000042004400000005004300000031004100000019004100000036004000000021004000000001003f0000001a003c00000008003c0000001f003b00000032003a0000001b003a0000001200380000002a00370000001000360000000600340000002500330000001700310000001500300000001e002d00000008002d00000020002c00000014002b00000023002a0000000b002a0000001700290000000700280000001c00270000000800240000001f00230000001a00220000000e00220000000c002000000018001f0000000a001f00000018001d00000015001d00000017001b00000003001b0000000d001a0000000b001a0000000e00190000000400190000000f00180000001000160000001300150000000000150000001000130000000b00120000000700110000000500110000000200100000000a000f0000000c000e00000007000d00000007000a0000000300090000000400080000000000080000000100050000001a00420001000600250000001600180000000a00160000000600150000000e00130000000100040000001d003500010024002f00010022002900010027002800010006002000010009001b00010000000300010015002e00000018002100000001001e00000014001a0000000c00190000000d00160000000f001400000008001400000010001200000002000f00000002000b0000000a00180000000800170000000c001000000012001600010013001c00000011001700000000001000000005000f00000009000e00000008000a0000000400070000000b001200010010001900000000001100000001001100000006000d0001000100150000000e000f00000002000400000005000700000006000c00000009000b0000000c000d00010002000f00010008000a00010011001200010000000400000007001400000005000e0000000900130001000100030000 ;
localparam YMAP = 1280'h000100ca000100be000000a6000100ba000000b4000000b7000000c2000100ae000000c7000000c1000000c5000100a8000100af000000b6000000ac000100b2000000a9000100a5000100bf000000b0000000b3000100bd000100b1000000bb000000c6000100a7000100c0000100aa000100b5000000c8000000ad00000084000000b8000000c4000000c3000000c9000000ab000100bc000100b90001007d;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 120'b010000001000100000001000000010001011010000000000000110000000000010010010111000100011000100011101000000100000000000000010 ;
localparam WNNZ = 120'b010000101000100000001000101010011011010000100010010110000000000010010010111001100011001100011101000000100001010000001010;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
wire [SUM_BITS-1:0] scorarr [CLASS_CNT-1:0];
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;

generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam adsub = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(adsub)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] <= 0;
end
endgenerate

function [7:0] zerocnt(input integer k);
    integer i,j;
    reg [HIDDEN_CNT-1:0] neur1;
    begin
        i = 0;
        neur1 = WNNZ[k*HIDDEN_CNT+:HIDDEN_CNT];
        for(j=0;j<HIDDEN_CNT;j=j+1)
            i = i + !(neur1[j]);
        zerocnt = i;
    end
endfunction

function [7:0] minzc(input integer k);
    integer i,j,h;
    begin
        i = HIDDEN_CNT;
        for(j=0;j<CLASS_CNT;j=j+1) begin
            h = zerocnt(j);
            if(h<i)
                i = h;
        end
        minzc = i;
    end
endfunction

localparam MINZC = minzc(0);

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    localparam Wuse = WNNZ[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wuse[j]) begin
            if(Wneur[j])
                tmpscore = tmpscore + hidden[j];
            else 
                tmpscore = tmpscore + hidden_n[j];
        end
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = 2*tmpscore + zerocnt(i) - MINZC;
    /* assign scorarr[i] = 2*tmpscore + zerocnt(i) - MINZC; */
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
