













module Har_bnn1_bnnroperm #(

parameter FEAT_CNT = 12,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 480'b000100000111011001111010001100000101000011110011000100101111101001101010000110110111001011101011000110000001100111001110111011101000111011111000101110101101011010001100000011000000101011110010000110010101111000010110111001100001111000111100100110000101011000001101000000100100101000111100110100000001110101000100110101010101111000110001001100101101100111100110010111110100001110000010100100000001110001110010001101001001111001110001010011011001110000111111010011110101101000111001 ;
  localparam Weights1 = 240'b100001111010000010011010111010111110101010100110101011111000010110111011100011101000011011100010001110101010111111001110000001100111111100010111101110100010010100000100001111010101100011111110010100110100000000010011010101001011101001100110 ;

  romesh_seq #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
