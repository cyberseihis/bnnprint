













module winewhite_bnn1_bnnroperm #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 440'b10011010110111110111110001111011000011001000001110101110110100011100111010010011110101101010111100010100111001011001111110110011110011100001000110000011000001011111111001011100100101000101111011100110010100010101101111010010011001100100010011001101100111101111111010001010101100011100110001110101010011001000110010010010101111001100110000101010100101111000010010100001011011000101010001001100110011000101001000000100110001000010011111010110 ;
  localparam Weights1 = 280'b0011101110100001100011000101000000111111011110111110010111010101010101100110101101111010111011011101010101010111010100110101100111100101010101000001011100000001011110111110010101010101010101110100001101111111101001011010110101010111010000111011101011110100110001010101001101000000 ;

  romesh_seq #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
