












module gasId_bnn1_bnndirect #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 5120'b00000110110011000100101101011001110011111100100010110010000010110100001101100101100110010111001101110000001110000110001011110110100011011101000001000111010100111111010010001101100110000000001001010110101010000000110111000010010101100100100110101010100010010001110000010110100011001110000100011010100001101001111010110101101001000110100011001001100000001010001110100001101011100001100110010110110101100101100011110110101000001100111111101111011101000000110100011000000110100001101011100100100011011001100000000011010111101010010110001101111011000111011011101100111100000000100110111100000101011001100010111001110110011100100100011111011111001101001011000011100000001011010000111101110101011100001100011110110110010001101100100011000001110010111000100100100111011111010010100101110110000000001001011011011001001010111011010010011000100101101101010101011001001011001011100010001110110001010001100011011101110000100100100011010101110111000010000010110010111011101100111100100001001100011000101111110001111100101110111000001001101010111011000100101000000001001001110011000011000010010011110100101011011001100000000010010110110101010010101111111111100110001001010011010000001110010000111110011000100101101011010110010100100111001100111011000010111101101111100000001000110110001110111011010101010001110101001011110010011100010110100101010101110001101010100110011010011111011010100010110100001010000100001101110001100000111101110111000111000001000011110000100011011101110100001011101100101010110010000000011101011101111110101110101000101101100001111100000011110110111000010011100010101100100111011111101010011111010110000001001101010010110100010000111001101110000110011111001001110001101110110110001101001001110011110000101100111010110000000001000010010000011010001010111001000000100110011000000100110100111010111000110010010110010110010111111011001011101000001001010111000001010110101110101100110011100010001000100111111110111110101001101100111101111011111010100110011000111111010001001111000011010001000001001111011110011111011011110101001101110001101001101010011100000001000010011100010111110010101111110000100110000001010001011110001010111011001000110010100101000101110100101011111111001011110010010100010111100010101101100000001110011001011101011111101001111111000110011000001101110001101101101101101000111111100000010110101110100111011100011001101001111111111000001010111011110011000000110001100111100100111010101011101100000011100100010100010110100010111110100000001110010001110101001101100010111001100110111111000001000100101011101011111100000011000100010101010000011100000110111000001111110011101100110100000101111110000000010101111010011010000011110110010011000101110011001010000110010010101111100101101001101101011000111001000010101110111000000110110001001001100110001011101001101010000011000101110001011011101010100111100111100011111001000000011011100011100111010101111010011001011010100101001011010010111011000010000011110010000110110111010101100111100011110100001010100001011011101001100001001111100100101010011101000001000000010110101100010010001101011111000001001101001111110001000100100000010000110110101110010000111101111011110111010111100000100111111010100110100000101011101100110111001111001011100010010010110111100110110001111001101010001001111111010100111101010111000010101000101101011011000001011010110100101111100101001000101100000111011011101011000100101001011101100001000010010110110100010001100110101001110110100010010001111101001011101001101111100100001100111101010101011100001011111000010000001010010101100111011001111001110000110101001111100111011011010111011111011100011011010011001111010111000010101010001101111001101001101110000010011011111110111110101001111001001010110111011000010000100101101101000100011001101110011111111010001110011011101110011111111000001010111110100001000010010101000110110010111010101011100000111110110110001001000101101000100000000001000111001010010010001000011110100011011000101110101100001111101100000011101001011100101011001001101011100000011110111011010001001111001111010001111110001110100010010101000000111111000011111010111011111100010110010111110100011111010011100100001101111000001010100101101010101111111111111111110111011101010101011101101100101011000010100110011101000001001100110101001011100101011010001101000001111011011001001011011101000100001000110011011010100011110010010001000100000111000011101100010101010101011111110001111110111110100010100100100100111101000111111110111001001001111100011101101101000011101011101100010011111111000010010110100101010000110111100001100011000011110111001011110110110000000010111101110101101110010010000011101111111000110010011100011110110101001010111011111001100111111101001001000100101011101011100000000011110100101101011010101110011010100000011000001011111101001110111011101011001000110001101111110100101011001111001111010011001001100011000100011011101100001001011000100101100100000011110100001100011001011100000011001110110010101111110101010110000010100100010010001010101111100001001110000011010001101010111010111110000101110011001101001001000011111111110101100010000010010100110011100010101110101000101110011001110101 ;
  localparam Weights1 = 240'b001101100010110011101111111110000101100100111011101110001100100011010110111110010011010000101000111011101111100011011101110101110110000001111111010010111010101110110110000010000111110101011111100011100111010010101100110110001100101001011011 ;

  seq_bnn #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
