`timescale 1us/1ns





module tbHar_tnn1_tnnseq #(

parameter FEAT_CNT = 12,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000




)();
  reg [FEAT_BITS*FEAT_CNT-1:0] data;
  wire [FEAT_BITS*FEAT_CNT-1:0] testcases [TEST_CNT-1:0];
  reg rst;
  reg clk;
  parameter Nsperiod=50000;
  localparam period=Nsperiod/500;
  localparam halfT=period/2;


assign testcases[0] = 48'h121a8941189b;
assign testcases[1] = 48'h011a7810079b;
assign testcases[2] = 48'h000a8800079b;
assign testcases[3] = 48'h000a8800079b;
assign testcases[4] = 48'h00098800079b;
assign testcases[5] = 48'h00098800079b;
assign testcases[6] = 48'h00099800079b;
assign testcases[7] = 48'h00098800079b;
assign testcases[8] = 48'h00098800079b;
assign testcases[9] = 48'h00098800079b;
assign testcases[10] = 48'h00098800079b;
assign testcases[11] = 48'h00098800079b;
assign testcases[12] = 48'h00098800079b;
assign testcases[13] = 48'h00098800079b;
assign testcases[14] = 48'h00099800079b;
assign testcases[15] = 48'h11299700079b;
assign testcases[16] = 48'h00088821179b;
assign testcases[17] = 48'h00098811079b;
assign testcases[18] = 48'h00098800079b;
assign testcases[19] = 48'h101a8801079b;
assign testcases[20] = 48'h101a8811078b;
assign testcases[21] = 48'h11199811079b;
assign testcases[22] = 48'h3219981118ab;
assign testcases[23] = 48'h3109881108ab;
assign testcases[24] = 48'h00098800079b;
assign testcases[25] = 48'h00098800079b;
assign testcases[26] = 48'h00098800079b;
assign testcases[27] = 48'h00098800079b;
assign testcases[28] = 48'h00098800079b;
assign testcases[29] = 48'h00098800079b;
assign testcases[30] = 48'h00098800079b;
assign testcases[31] = 48'h100a8811079b;
assign testcases[32] = 48'h000a9800079b;
assign testcases[33] = 48'h00098800079b;
assign testcases[34] = 48'h00098800079b;
assign testcases[35] = 48'h00098800079b;
assign testcases[36] = 48'h00098800079b;
assign testcases[37] = 48'h00098800079b;
assign testcases[38] = 48'h00098800079b;
assign testcases[39] = 48'h00098800079b;
assign testcases[40] = 48'h00098800079b;
assign testcases[41] = 48'h00098800079b;
assign testcases[42] = 48'h00098800079b;
assign testcases[43] = 48'h00098800079b;
assign testcases[44] = 48'h2115a62116ab;
assign testcases[45] = 48'h20179711079b;
assign testcases[46] = 48'h10099700079b;
assign testcases[47] = 48'h00098800079b;
assign testcases[48] = 48'h00098800079b;
assign testcases[49] = 48'h100a8800079b;
assign testcases[50] = 48'h000a8801079b;
assign testcases[51] = 48'h00098800078b;
assign testcases[52] = 48'h00098800079b;
assign testcases[53] = 48'h00099800079b;
assign testcases[54] = 48'h00098800079b;
assign testcases[55] = 48'h111b6800179a;
assign testcases[56] = 48'h110a7800079b;
assign testcases[57] = 48'h00098800079b;
assign testcases[58] = 48'h00098800079b;
assign testcases[59] = 48'h00099800079b;
assign testcases[60] = 48'h00099800079b;
assign testcases[61] = 48'h00099800079b;
assign testcases[62] = 48'h00098800079b;
assign testcases[63] = 48'h00098800079b;
assign testcases[64] = 48'h00098800079b;
assign testcases[65] = 48'h00098800079b;
assign testcases[66] = 48'h201e6911279c;
assign testcases[67] = 48'h211b6800179c;
assign testcases[68] = 48'h100a7800079b;
assign testcases[69] = 48'h10098800079b;
assign testcases[70] = 48'h00098800079b;
assign testcases[71] = 48'h00098800079b;
assign testcases[72] = 48'h00099800079b;
assign testcases[73] = 48'h00098800079b;
assign testcases[74] = 48'h00098800079b;
assign testcases[75] = 48'h00099800079b;
assign testcases[76] = 48'h00098800079b;
assign testcases[77] = 48'h00098800079c;
assign testcases[78] = 48'h00099800079b;
assign testcases[79] = 48'h6549b667679a;
assign testcases[80] = 48'h654a9767789b;
assign testcases[81] = 48'h55498878679c;
assign testcases[82] = 48'h55498878579b;
assign testcases[83] = 48'h55498877579b;
assign testcases[84] = 48'h55498866679a;
assign testcases[85] = 48'h6549886667ab;
assign testcases[86] = 48'h64498867679c;
assign testcases[87] = 48'h65499877679c;
assign testcases[88] = 48'h55599767579c;
assign testcases[89] = 48'h655a9867679a;
assign testcases[90] = 48'h75599877689a;
assign testcases[91] = 48'h65599877679c;
assign testcases[92] = 48'h55598867679b;
assign testcases[93] = 48'h654a786667aa;
assign testcases[94] = 48'h5549c566679b;
assign testcases[95] = 48'h5549a677778c;
assign testcases[96] = 48'h65599767779a;
assign testcases[97] = 48'h555a886768ab;
assign testcases[98] = 48'h55498867679c;
assign testcases[99] = 48'h55498867678b;
assign testcases[100] = 48'h5559886767ab;
assign testcases[101] = 48'h5549886767ab;
assign testcases[102] = 48'h65598867679c;
assign testcases[103] = 48'h65599867778b;
assign testcases[104] = 48'h554a9767679a;
assign testcases[105] = 48'h5549887768ab;
assign testcases[106] = 48'h65499878678c;
assign testcases[107] = 48'h55499868678b;
assign testcases[108] = 48'h55498877579b;
assign testcases[109] = 48'h64499788978c;
assign testcases[110] = 48'h65399778a69c;
assign testcases[111] = 48'h7479b69998ab;
assign testcases[112] = 48'h7469b5999899;
assign testcases[113] = 48'h755a78799798;
assign testcases[114] = 48'h7689a78aa79c;
assign testcases[115] = 48'h7789979ab7ab;
assign testcases[116] = 48'h86595baab78b;
assign testcases[117] = 48'h86496b99a78d;
assign testcases[118] = 48'h664b96a9a69b;
assign testcases[119] = 48'h764a97b8b69c;
assign testcases[120] = 48'h878bd4dab69d;
assign testcases[121] = 48'h87aa96cbb69a;
assign testcases[122] = 48'h86aa87bab7aa;
assign testcases[123] = 48'h879a97caa79b;
assign testcases[124] = 48'h76677bcac78b;
assign testcases[125] = 48'h86676acad89b;
assign testcases[126] = 48'h857fb4eae78b;
assign testcases[127] = 48'h868fc3d8b7ab;
assign testcases[128] = 48'ha79db5d8a79b;
assign testcases[129] = 48'h977a98dab8ab;
assign testcases[130] = 48'h979a97ebc69d;
assign testcases[131] = 48'h96a769e9c78a;
assign testcases[132] = 48'h76655cdab79a;
assign testcases[133] = 48'h9649b4b9739b;
assign testcases[134] = 48'ha749b689748a;
assign testcases[135] = 48'ha6588988779a;
assign testcases[136] = 48'h95765b8867ab;
assign testcases[137] = 48'h967979a9769b;
assign testcases[138] = 48'hc7689888769a;
assign testcases[139] = 48'hc6788978779a;
assign testcases[140] = 48'ha66ca6b885ab;
assign testcases[141] = 48'ha73bb5b875ab;
assign testcases[142] = 48'ha65b94c97398;
assign testcases[143] = 48'hb67aa7d873ba;
assign testcases[144] = 48'hd6779ab8769b;
assign testcases[145] = 48'hc5757ba9779b;
assign testcases[146] = 48'hb58a99ba779a;
assign testcases[147] = 48'he67889ba86ab;
assign testcases[148] = 48'hf78988c977ab;
assign testcases[149] = 48'hb67fb5c87799;
assign testcases[150] = 48'hb56eb5c97568;
assign testcases[151] = 48'ha47aa7d8769b;
assign testcases[152] = 48'hf5747ab9679b;
assign testcases[153] = 48'hf5757ac9679b;
assign testcases[154] = 48'hb47a98c8669b;
assign testcases[155] = 48'hd68889d9679a;
assign testcases[156] = 48'hd78c97e9789b;
assign testcases[157] = 48'ha67fa5e9778b;
assign testcases[158] = 48'h11198941188a;
assign testcases[159] = 48'h001a8801069b;
assign testcases[160] = 48'h000a8800069b;
assign testcases[161] = 48'h000a8810079b;
assign testcases[162] = 48'h00099800079b;
assign testcases[163] = 48'h00099800079b;
assign testcases[164] = 48'h00098800079b;
assign testcases[165] = 48'h00098800079b;
assign testcases[166] = 48'h00098800079b;
assign testcases[167] = 48'h00098800079b;
assign testcases[168] = 48'h00098800079b;
assign testcases[169] = 48'h1008983108ac;
assign testcases[170] = 48'h00098800069b;
assign testcases[171] = 48'h00098800079b;
assign testcases[172] = 48'h00098800079b;
assign testcases[173] = 48'h00098800079b;
assign testcases[174] = 48'h00098800079b;
assign testcases[175] = 48'h00098800079b;
assign testcases[176] = 48'h00098800079b;
assign testcases[177] = 48'h00098800079b;
assign testcases[178] = 48'h00098800079b;
assign testcases[179] = 48'h00098800079b;
assign testcases[180] = 48'h10099800079b;
assign testcases[181] = 48'h110a882208cb;
assign testcases[182] = 48'h100a881108aa;
assign testcases[183] = 48'h000a8800079b;
assign testcases[184] = 48'h000a8800079b;
assign testcases[185] = 48'h00098800079b;
assign testcases[186] = 48'h00098800079b;
assign testcases[187] = 48'h00098800079b;
assign testcases[188] = 48'h00098800079b;
assign testcases[189] = 48'h00098800079b;
assign testcases[190] = 48'h00099800079b;
assign testcases[191] = 48'h00098800079b;
assign testcases[192] = 48'h1102b654235d;
assign testcases[193] = 48'h2014a710079b;
assign testcases[194] = 48'h2006a700079b;
assign testcases[195] = 48'h10089800079b;
assign testcases[196] = 48'h00098800079b;
assign testcases[197] = 48'h000a8800079b;
assign testcases[198] = 48'h00098800079b;
assign testcases[199] = 48'h00098800079b;
assign testcases[200] = 48'h00098800079b;
assign testcases[201] = 48'h00098800079b;
assign testcases[202] = 48'h00098800079b;
assign testcases[203] = 48'h210f7811269b;
assign testcases[204] = 48'h200d7800179b;
assign testcases[205] = 48'h100b8800079a;
assign testcases[206] = 48'h00098800079b;
assign testcases[207] = 48'h00098800079b;
assign testcases[208] = 48'h00099800079b;
assign testcases[209] = 48'h00099800079b;
assign testcases[210] = 48'h00098800079b;
assign testcases[211] = 48'h00098800079b;
assign testcases[212] = 48'h00098800079b;
assign testcases[213] = 48'h00098800079b;
assign testcases[214] = 48'h211d7911179b;
assign testcases[215] = 48'h100b7800079b;
assign testcases[216] = 48'h00098800079b;
assign testcases[217] = 48'h00098800079b;
assign testcases[218] = 48'h00099800079b;
assign testcases[219] = 48'h00098800079b;
assign testcases[220] = 48'h00098800079b;
assign testcases[221] = 48'h00099800079b;
assign testcases[222] = 48'h00098800079b;
assign testcases[223] = 48'h00098800079b;
assign testcases[224] = 48'h00098800079b;
assign testcases[225] = 48'h00098800079b;
assign testcases[226] = 48'h00098800079b;
assign testcases[227] = 48'h5558c567687b;
assign testcases[228] = 48'h66699668779a;
assign testcases[229] = 48'h66598868879b;
assign testcases[230] = 48'h655a8867679b;
assign testcases[231] = 48'h554a885857ab;
assign testcases[232] = 48'h64498868679b;
assign testcases[233] = 48'h64599868678c;
assign testcases[234] = 48'h55599867679a;
assign testcases[235] = 48'h65598867689b;
assign testcases[236] = 48'h65598868679c;
assign testcases[237] = 48'h65598868769a;
assign testcases[238] = 48'h6559885867aa;
assign testcases[239] = 48'h64599867679c;
assign testcases[240] = 48'h64598867579c;
assign testcases[241] = 48'h54599857579b;
assign testcases[242] = 48'h7668b568779c;
assign testcases[243] = 48'h76699678879b;
assign testcases[244] = 48'h77699779779b;
assign testcases[245] = 48'h666a8869679b;
assign testcases[246] = 48'h655a886767aa;
assign testcases[247] = 48'h65598868779c;
assign testcases[248] = 48'h65699768779b;
assign testcases[249] = 48'h65698868779b;
assign testcases[250] = 48'h6659887a779c;
assign testcases[251] = 48'h66598879779a;
assign testcases[252] = 48'h6649886767ab;
assign testcases[253] = 48'h66599867679c;
assign testcases[254] = 48'h66599867679b;
assign testcases[255] = 48'h55498856679b;
assign testcases[256] = 48'h955998a9c69c;
assign testcases[257] = 48'h86598899c899;
assign testcases[258] = 48'h7688b57ab79b;
assign testcases[259] = 48'h9788b58bb79b;
assign testcases[260] = 48'ha788978bc79b;
assign testcases[261] = 48'h8779976aa6ac;
assign testcases[262] = 48'h887b6a8cb78b;
assign testcases[263] = 48'h887b6b8cc68b;
assign testcases[264] = 48'h7568e38ae88b;
assign testcases[265] = 48'h8687d38cd89b;
assign testcases[266] = 48'h8687c39dd6ab;
assign testcases[267] = 48'h8879889cd79b;
assign testcases[268] = 48'h8899979bd69b;
assign testcases[269] = 48'h88b9989ce78b;
assign testcases[270] = 48'h878a5c8cd89a;
assign testcases[271] = 48'h9778d48ac78a;
assign testcases[272] = 48'h9868b589c89d;
assign testcases[273] = 48'h9997d39ac69b;
assign testcases[274] = 48'h88b996aac789;
assign testcases[275] = 48'h7799a78ac89a;
assign testcases[276] = 48'h88b9988cd79d;
assign testcases[277] = 48'h977b5c8cd7ab;
assign testcases[278] = 48'h967b7a7bd79b;
assign testcases[279] = 48'h7549d48a964a;
assign testcases[280] = 48'h6648b68a978c;
assign testcases[281] = 48'h77885b8987ab;
assign testcases[282] = 48'h87995b89879b;
assign testcases[283] = 48'h75499789868b;
assign testcases[284] = 48'h75597988779b;
assign testcases[285] = 48'h666aa798779b;
assign testcases[286] = 48'h6639d57887aa;
assign testcases[287] = 48'h6558b599848a;
assign testcases[288] = 48'h7559978a978b;
assign testcases[289] = 48'h75795a99979c;
assign testcases[290] = 48'h76695b89879b;
assign testcases[291] = 48'h7649888a988b;
assign testcases[292] = 48'h8679798a87ab;
assign testcases[293] = 48'h7789978986aa;
assign testcases[294] = 48'h7639b57997aa;
assign testcases[295] = 48'h6658c599948c;
assign testcases[296] = 48'h76688889979c;
assign testcases[297] = 48'h76596a8a889b;
assign testcases[298] = 48'h6769998a97ab;
assign testcases[299] = 48'h6769798987ab;
assign testcases[300] = 48'h768a8878879b;
assign testcases[301] = 48'h654ad478889a;
assign testcases[302] = 48'h332aaa741daa;
assign testcases[303] = 48'h314a8842167b;
assign testcases[304] = 48'h11298722069b;
assign testcases[305] = 48'h1119872008ab;
assign testcases[306] = 48'h1129872108ab;
assign testcases[307] = 48'h21398811079b;
assign testcases[308] = 48'h21199811079b;
assign testcases[309] = 48'h1119881107ab;
assign testcases[310] = 48'h00098800079b;
assign testcases[311] = 48'h00098800079b;
assign testcases[312] = 48'h00098800079b;
assign testcases[313] = 48'h00098800079b;
assign testcases[314] = 48'h00198800079b;
assign testcases[315] = 48'h00098800079b;
assign testcases[316] = 48'h00198810079b;
assign testcases[317] = 48'h10399710079b;
assign testcases[318] = 48'h1018882417cc;
assign testcases[319] = 48'h10098810069b;
assign testcases[320] = 48'h000a8800079b;
assign testcases[321] = 48'h000a9800079b;
assign testcases[322] = 48'h10099800079b;
assign testcases[323] = 48'h00098801079b;
assign testcases[324] = 48'h10198801079b;
assign testcases[325] = 48'h10198801079b;
assign testcases[326] = 48'h00098801079b;
assign testcases[327] = 48'h00098800079b;
assign testcases[328] = 48'h10198800079b;
assign testcases[329] = 48'h11498731059b;
assign testcases[330] = 48'h100b881317ba;
assign testcases[331] = 48'h100b8800079b;
assign testcases[332] = 48'h000a8800079b;
assign testcases[333] = 48'h000a8800079b;
assign testcases[334] = 48'h00098800079b;
assign testcases[335] = 48'h00098800079b;
assign testcases[336] = 48'h00098800079b;
assign testcases[337] = 48'h00098800079b;
assign testcases[338] = 48'h00099800079b;
assign testcases[339] = 48'h00098800079b;
assign testcases[340] = 48'h00098800079b;
assign testcases[341] = 48'h100a8800079b;
assign testcases[342] = 48'h1016861107ab;
assign testcases[343] = 48'h1018870007ab;
assign testcases[344] = 48'h11098701079b;
assign testcases[345] = 48'h100a8801079b;
assign testcases[346] = 48'h000a8801079b;
assign testcases[347] = 48'h00098800079b;
assign testcases[348] = 48'h00098800079b;
assign testcases[349] = 48'h00099800079b;
assign testcases[350] = 48'h10099801079b;
assign testcases[351] = 48'h1009880107ab;
assign testcases[352] = 48'h00098801079b;
assign testcases[353] = 48'h110a8801079b;
assign testcases[354] = 48'h211f792347a8;
assign testcases[355] = 48'h111c7811179b;
assign testcases[356] = 48'h100b8800079a;
assign testcases[357] = 48'h000a8800079b;
assign testcases[358] = 48'h00098800079b;
assign testcases[359] = 48'h00098800079b;
assign testcases[360] = 48'h00098800079b;
assign testcases[361] = 48'h00099800079b;
assign testcases[362] = 48'h00098800079b;
assign testcases[363] = 48'h00098800079b;
assign testcases[364] = 48'h00098800079b;
assign testcases[365] = 48'h00098800079b;
assign testcases[366] = 48'h00098800079b;
assign testcases[367] = 48'h00098800079b;
assign testcases[368] = 48'h00099800079b;
assign testcases[369] = 48'h11098800079b;
assign testcases[370] = 48'h212e7923269c;
assign testcases[371] = 48'h212c792216ac;
assign testcases[372] = 48'h100a8810079b;
assign testcases[373] = 48'h00098800079b;
assign testcases[374] = 48'h00098800079b;
assign testcases[375] = 48'h00099800079b;
assign testcases[376] = 48'h00099800079b;
assign testcases[377] = 48'h00098800079b;
assign testcases[378] = 48'h00098800079b;
assign testcases[379] = 48'h00098800079b;
assign testcases[380] = 48'h00098800079b;
assign testcases[381] = 48'h00098800079b;
assign testcases[382] = 48'h00098800079b;
assign testcases[383] = 48'h00098800079b;
assign testcases[384] = 48'h4348965657bb;
assign testcases[385] = 48'h44599747679b;
assign testcases[386] = 48'h445a9756679b;
assign testcases[387] = 48'h34498856679b;
assign testcases[388] = 48'h34598847679b;
assign testcases[389] = 48'h4459984767ac;
assign testcases[390] = 48'h54599857679b;
assign testcases[391] = 48'h44598857678b;
assign testcases[392] = 48'h44598858669b;
assign testcases[393] = 48'h43598847579b;
assign testcases[394] = 48'h43499847679c;
assign testcases[395] = 48'h433a985668ab;
assign testcases[396] = 48'h33499766679b;
assign testcases[397] = 48'h34598857578b;
assign testcases[398] = 48'h4459885657ab;
assign testcases[399] = 48'h4359884757ac;
assign testcases[400] = 48'h54598b67668b;
assign testcases[401] = 48'h53598957679b;
assign testcases[402] = 48'h5359974867ab;
assign testcases[403] = 48'h445a9757679b;
assign testcases[404] = 48'h53598857678b;
assign testcases[405] = 48'h5469885867ab;
assign testcases[406] = 48'h4469885867ac;
assign testcases[407] = 48'h54599758679b;
assign testcases[408] = 48'h44698857678b;
assign testcases[409] = 48'h44598858679b;
assign testcases[410] = 48'h4459885867ac;
assign testcases[411] = 48'h44599757679b;
assign testcases[412] = 48'h43599856679b;
assign testcases[413] = 48'h44498857679b;
assign testcases[414] = 48'h4459885867ab;
assign testcases[415] = 48'h53598855a8ac;
assign testcases[416] = 48'h5359875597aa;
assign testcases[417] = 48'h53889466a79c;
assign testcases[418] = 48'h534a8b45b8aa;
assign testcases[419] = 48'h534a8a45c79b;
assign testcases[420] = 48'h5348a55488aa;
assign testcases[421] = 48'h5349975498ab;
assign testcases[422] = 48'h53499655979c;
assign testcases[423] = 48'h53889457878c;
assign testcases[424] = 48'h63a98657879b;
assign testcases[425] = 48'h537998658899;
assign testcases[426] = 48'h64899776879a;
assign testcases[427] = 48'h645a8a65969a;
assign testcases[428] = 48'h534a7a55b79b;
assign testcases[429] = 48'h53aa9666c69e;
assign testcases[430] = 48'h5458a565b8ac;
assign testcases[431] = 48'h53598655b8aa;
assign testcases[432] = 48'h63789456a79a;
assign testcases[433] = 48'h63989656978a;
assign testcases[434] = 48'h54899765a7ab;
assign testcases[435] = 48'h54999766979b;
assign testcases[436] = 48'h636a6b47b79c;
assign testcases[437] = 48'h635b8b56c6ac;
assign testcases[438] = 48'h84387878857c;
assign testcases[439] = 48'h8449876687aa;
assign testcases[440] = 48'h844989668899;
assign testcases[441] = 48'h645b8b77889b;
assign testcases[442] = 48'h746a9977769b;
assign testcases[443] = 48'h94489657869c;
assign testcases[444] = 48'h94797967779b;
assign testcases[445] = 48'h94697967779a;
assign testcases[446] = 48'h9449a667878c;
assign testcases[447] = 48'h744aa667879c;
assign testcases[448] = 48'h745aa66677aa;
assign testcases[449] = 48'h845a8967976a;
assign testcases[450] = 48'h74598866979b;
assign testcases[451] = 48'h656a8a77889c;
assign testcases[452] = 48'h656b7b68879c;
assign testcases[453] = 48'h75798867869b;
assign testcases[454] = 48'h856a8978979b;
assign testcases[455] = 48'h85699878979b;
assign testcases[456] = 48'h8558a578978b;
assign testcases[457] = 48'h85699668979b;
assign testcases[458] = 48'h856a9b79a66c;
assign testcases[459] = 48'h75699967a88c;
assign testcases[460] = 48'h856a6b77879b;
assign testcases[461] = 48'h85897a78979b;
assign testcases[462] = 48'h85799768979b;
assign testcases[463] = 48'h857a7988989b;
assign testcases[464] = 48'h75899687969b;
assign testcases[465] = 48'h7569b477969b;
assign testcases[466] = 48'h6414f8573efc;
assign testcases[467] = 48'h3219b862199a;
assign testcases[468] = 48'h21299811068b;
assign testcases[469] = 48'h21198721069b;
assign testcases[470] = 48'h201a8812079b;
assign testcases[471] = 48'h101a8811079b;
assign testcases[472] = 48'h10198800079b;
assign testcases[473] = 48'h10198701079b;
assign testcases[474] = 48'h10199801079b;
assign testcases[475] = 48'h10199811079b;
assign testcases[476] = 48'h10199811089b;
assign testcases[477] = 48'h10198811079b;
assign testcases[478] = 48'h10198811079b;
assign testcases[479] = 48'h00098810079b;
assign testcases[480] = 48'h00098810079b;
assign testcases[481] = 48'h111a8812078b;
assign testcases[482] = 48'h2127882718ed;
assign testcases[483] = 48'h10188812078b;
assign testcases[484] = 48'h10198711079b;
assign testcases[485] = 48'h10298801079b;
assign testcases[486] = 48'h1029980207ab;
assign testcases[487] = 48'h101a871207ab;
assign testcases[488] = 48'h101a8801078b;
assign testcases[489] = 48'h10198811079b;
assign testcases[490] = 48'h1009880106ab;
assign testcases[491] = 48'h100a9811079b;
assign testcases[492] = 48'h00099800088b;
assign testcases[493] = 48'h10198811079b;
assign testcases[494] = 48'h110d881917d8;
assign testcases[495] = 48'h100c8801078b;
assign testcases[496] = 48'h100b8800079b;
assign testcases[497] = 48'h100a8800079b;
assign testcases[498] = 48'h00098800079b;
assign testcases[499] = 48'h10099801079b;
assign testcases[500] = 48'h10099811079b;
assign testcases[501] = 48'h11098801079b;
assign testcases[502] = 48'h11098811079b;
assign testcases[503] = 48'h01098800069b;
assign testcases[504] = 48'h00098800079b;
assign testcases[505] = 48'h00099800079b;
assign testcases[506] = 48'h00098800079b;
assign testcases[507] = 48'h00098800079b;
assign testcases[508] = 48'h513575951adb;
assign testcases[509] = 48'h21187611058b;
assign testcases[510] = 48'h10198701078b;
assign testcases[511] = 48'h10198801079b;
assign testcases[512] = 48'h10098801079b;
assign testcases[513] = 48'h1009980107ab;
assign testcases[514] = 48'h11199811079b;
assign testcases[515] = 48'h1119981108ab;
assign testcases[516] = 48'h1109881107bb;
assign testcases[517] = 48'h320a8823178b;
assign testcases[518] = 48'h320a9823188b;
assign testcases[519] = 48'h12198821079b;
assign testcases[520] = 48'h211f992468b4;
assign testcases[521] = 48'h111d9901179c;
assign testcases[522] = 48'h100b8800079b;
assign testcases[523] = 48'h100a8801079b;
assign testcases[524] = 48'h11198811079b;
assign testcases[525] = 48'h10098811079b;
assign testcases[526] = 48'h00098800079b;
assign testcases[527] = 48'h00098800079b;
assign testcases[528] = 48'h00099800079b;
assign testcases[529] = 48'h00098800079b;
assign testcases[530] = 48'h00098800079b;
assign testcases[531] = 48'h00099801079b;
assign testcases[532] = 48'h111f89234898;
assign testcases[533] = 48'h211d8811179c;
assign testcases[534] = 48'h100b8800079b;
assign testcases[535] = 48'h100a8800079b;
assign testcases[536] = 48'h00098800079b;
assign testcases[537] = 48'h00098800079b;
assign testcases[538] = 48'h00098800079b;
assign testcases[539] = 48'h00098800079b;
assign testcases[540] = 48'h00099800079b;
assign testcases[541] = 48'h00098800079b;
assign testcases[542] = 48'h00098800079b;
assign testcases[543] = 48'h00099800079b;
assign testcases[544] = 48'h43488847669b;
assign testcases[545] = 48'h335a974767ab;
assign testcases[546] = 48'h34599747678b;
assign testcases[547] = 48'h34598848679b;
assign testcases[548] = 48'h3469884877ab;
assign testcases[549] = 48'h44699748679b;
assign testcases[550] = 48'h34698848679b;
assign testcases[551] = 48'h3469884867ab;
assign testcases[552] = 48'h33698848679c;
assign testcases[553] = 48'h34599747688b;
assign testcases[554] = 48'h34599848679b;
assign testcases[555] = 48'h34598848679b;
assign testcases[556] = 48'h34598848779b;
assign testcases[557] = 48'h34599747779b;
assign testcases[558] = 48'h44e8924756ab;
assign testcases[559] = 48'h445a8b48678b;
assign testcases[560] = 48'h346a894776ab;
assign testcases[561] = 48'h33699748779b;
assign testcases[562] = 48'h43698849779b;
assign testcases[563] = 48'h44698849779b;
assign testcases[564] = 48'h4469a748779b;
assign testcases[565] = 48'h34699848779a;
assign testcases[566] = 48'h33598849679b;
assign testcases[567] = 48'h34698848769b;
assign testcases[568] = 48'h34799748779b;
assign testcases[569] = 48'h34798848789a;
assign testcases[570] = 48'h34698849679b;
assign testcases[571] = 48'h34699839669c;
assign testcases[572] = 48'h3469974768ab;
assign testcases[573] = 48'h53588766c79c;
assign testcases[574] = 48'h43598766c8ac;
assign testcases[575] = 48'h63788468b78c;
assign testcases[576] = 48'h74998768b79a;
assign testcases[577] = 48'h548a9766a7aa;
assign testcases[578] = 48'h53998867b68a;
assign testcases[579] = 48'h535a8b66d79a;
assign testcases[580] = 48'h536a9956e6ac;
assign testcases[581] = 48'h63689666d7ab;
assign testcases[582] = 48'h5358a556c6ab;
assign testcases[583] = 48'h64979467b78b;
assign testcases[584] = 48'h73a88668c89d;
assign testcases[585] = 48'h63998768c79c;
assign testcases[586] = 48'h639a7958d789;
assign testcases[587] = 48'h536b7b67f6aa;
assign testcases[588] = 48'h53589566e7ac;
assign testcases[589] = 48'h5468a468d7ab;
assign testcases[590] = 48'h74a89478c78c;
assign testcases[591] = 48'h74a88667c79b;
assign testcases[592] = 48'h53898767c8a9;
assign testcases[593] = 48'h838a7a77d79c;
assign testcases[594] = 48'h847b8b69d59b;
assign testcases[595] = 48'h76598b88a66a;
assign testcases[596] = 48'h66598a87989b;
assign testcases[597] = 48'h666a6b8798ac;
assign testcases[598] = 48'h66798987979b;
assign testcases[599] = 48'h76698778978b;
assign testcases[600] = 48'h75797968978b;
assign testcases[601] = 48'h66889677969a;
assign testcases[602] = 48'h6669a477969a;
assign testcases[603] = 48'h756a8a78a76b;
assign testcases[604] = 48'h66598978a79c;
assign testcases[605] = 48'h765a7b68979c;
assign testcases[606] = 48'h75798a78979b;
assign testcases[607] = 48'h66598878989a;
assign testcases[608] = 48'h666a8978879b;
assign testcases[609] = 48'h5579b67896aa;
assign testcases[610] = 48'h6559a57897aa;
assign testcases[611] = 48'h657a8c79a64b;
assign testcases[612] = 48'h55798b78a79a;
assign testcases[613] = 48'h86696c7897aa;
assign testcases[614] = 48'h86898a78989b;
assign testcases[615] = 48'h657a988788ac;
assign testcases[616] = 48'h56698877978b;
assign testcases[617] = 48'h56599477978a;
assign testcases[618] = 48'h66789677969a;
assign testcases[619] = 48'h121a982118ab;
assign testcases[620] = 48'h101a8810079b;
assign testcases[621] = 48'h00099810079b;
assign testcases[622] = 48'h00098810079b;
assign testcases[623] = 48'h00098810079b;
assign testcases[624] = 48'h00098800079b;
assign testcases[625] = 48'h00098800079b;
assign testcases[626] = 48'h00099800079b;
assign testcases[627] = 48'h00098800079b;
assign testcases[628] = 48'h00098800079b;
assign testcases[629] = 48'h00198830089b;
assign testcases[630] = 48'h00198810079b;
assign testcases[631] = 48'h00098800079b;
assign testcases[632] = 48'h00098800079b;
assign testcases[633] = 48'h00098800079b;
assign testcases[634] = 48'h00098800079b;
assign testcases[635] = 48'h00098800079b;
assign testcases[636] = 48'h10399701079b;
assign testcases[637] = 48'h22498811168b;
assign testcases[638] = 48'h22298821169b;
assign testcases[639] = 48'h1119981108ab;
assign testcases[640] = 48'h1119982108ab;
assign testcases[641] = 48'h111a8822189a;
assign testcases[642] = 48'h000a8810079b;
assign testcases[643] = 48'h000a8800079b;
assign testcases[644] = 48'h00098800079b;
assign testcases[645] = 48'h00099800079b;
assign testcases[646] = 48'h00098800079b;
assign testcases[647] = 48'h00098800079b;
assign testcases[648] = 48'h00098800079b;
assign testcases[649] = 48'h00098800079b;
assign testcases[650] = 48'h00098800079b;
assign testcases[651] = 48'h00098800079b;
assign testcases[652] = 48'h1117e621189b;
assign testcases[653] = 48'h1119b710079b;
assign testcases[654] = 48'h01099710079b;
assign testcases[655] = 48'h00098800079b;
assign testcases[656] = 48'h00098810079b;
assign testcases[657] = 48'h01098811079b;
assign testcases[658] = 48'h00098811079b;
assign testcases[659] = 48'h1009881107ab;
assign testcases[660] = 48'h01099811079b;
assign testcases[661] = 48'h01098811079b;
assign testcases[662] = 48'h01098811079b;
assign testcases[663] = 48'h00099810079b;
assign testcases[664] = 48'h00098810079b;
assign testcases[665] = 48'h00098800079b;
assign testcases[666] = 48'h122c28438892;
assign testcases[667] = 48'h131b4821179c;
assign testcases[668] = 48'h121a6821179b;
assign testcases[669] = 48'h11198810179a;
assign testcases[670] = 48'h01099810179a;
assign testcases[671] = 48'h00098800179a;
assign testcases[672] = 48'h00098800079b;
assign testcases[673] = 48'h01098800079b;
assign testcases[674] = 48'h01098800079b;
assign testcases[675] = 48'h00098800079b;
assign testcases[676] = 48'h00098800079b;
assign testcases[677] = 48'h00098800079b;
assign testcases[678] = 48'h212c39131779;
assign testcases[679] = 48'h111b5911178a;
assign testcases[680] = 48'h110a7800079b;
assign testcases[681] = 48'h01098801079b;
assign testcases[682] = 48'h00099800079b;
assign testcases[683] = 48'h01198811179c;
assign testcases[684] = 48'h11199811179b;
assign testcases[685] = 48'h11199801079b;
assign testcases[686] = 48'h01199811179b;
assign testcases[687] = 48'h01199811179a;
assign testcases[688] = 48'h01098800179b;
assign testcases[689] = 48'h00098800079b;
assign testcases[690] = 48'h855aa8a7868b;
assign testcases[691] = 48'h856998a7889b;
assign testcases[692] = 48'h866889a787ab;
assign testcases[693] = 48'h956988a7979b;
assign testcases[694] = 48'h956a97a7979b;
assign testcases[695] = 48'h857998b7879b;
assign testcases[696] = 48'h857988a788ab;
assign testcases[697] = 48'h74598895779b;
assign testcases[698] = 48'h645a89a5679b;
assign testcases[699] = 48'h646987a6679b;
assign testcases[700] = 48'h6459879667aa;
assign testcases[701] = 48'h755998a6679c;
assign testcases[702] = 48'h745988a6779b;
assign testcases[703] = 48'h656ab3b6868a;
assign testcases[704] = 48'h746a94a6879b;
assign testcases[705] = 48'h84699797869b;
assign testcases[706] = 48'h8458889677ab;
assign testcases[707] = 48'h855988a6879b;
assign testcases[708] = 48'h856a98a7878b;
assign testcases[709] = 48'h867998a7879b;
assign testcases[710] = 48'h857989a887ab;
assign testcases[711] = 48'h856988a798ab;
assign testcases[712] = 48'h855a8797889b;
assign testcases[713] = 48'h84599796878b;
assign testcases[714] = 48'h85699897779a;
assign testcases[715] = 48'h7449899777ab;
assign testcases[716] = 48'h65499866b99c;
assign testcases[717] = 48'h65698666d79c;
assign testcases[718] = 48'h75999965d89c;
assign testcases[719] = 48'h86899675c59d;
assign testcases[720] = 48'h85799975b8a9;
assign testcases[721] = 48'h655a8b76c89b;
assign testcases[722] = 48'h76698876d68d;
assign testcases[723] = 48'h755cb066679a;
assign testcases[724] = 48'h845a9466668b;
assign testcases[725] = 48'h84488666659c;
assign testcases[726] = 48'h83489765468a;
assign testcases[727] = 48'h959a8a7667ab;
assign testcases[728] = 48'ha4898875668a;
assign testcases[729] = 48'ha4798976689c;
assign testcases[730] = 48'ha45a956568ac;
assign testcases[731] = 48'h945b9465679b;
assign testcases[732] = 48'h95c89a66669a;
assign testcases[733] = 48'h856aa376c8aa;
assign testcases[734] = 48'h765b8566c79b;
assign testcases[735] = 48'h986ba69acaab;
assign testcases[736] = 48'h989996aad88b;
assign testcases[737] = 48'ha8a888a8e79c;
assign testcases[738] = 48'h875a8b86e7aa;
assign testcases[739] = 48'ha46aa366757b;
assign testcases[740] = 48'hb47aa665767b;
assign testcases[741] = 48'hd5889a87679a;
assign testcases[742] = 48'hc679898777ab;
assign testcases[743] = 48'h9569986568ab;
assign testcases[744] = 48'ha5598a65679b;
assign testcases[745] = 48'hb57b8666768c;
assign testcases[746] = 48'ha56a9566778c;
assign testcases[747] = 48'h777aa476d9aa;
assign testcases[748] = 48'h667a8476e89d;
assign testcases[749] = 48'h66699387e68c;
assign testcases[750] = 48'h789887b8f69a;
assign testcases[751] = 48'h88aa97caf58b;
assign testcases[752] = 48'h8799a8aad9ab;
assign testcases[753] = 48'h86597c87eaba;
assign testcases[754] = 48'h785a7b76f78b;
assign testcases[755] = 48'hb46ab276658b;
assign testcases[756] = 48'hb468a366569a;
assign testcases[757] = 48'hb5968977679b;
assign testcases[758] = 48'hc5898a7777ac;
assign testcases[759] = 48'hc56a9967779b;
assign testcases[760] = 48'hc55a8977678a;
assign testcases[761] = 48'hb65b8677679b;
assign testcases[762] = 48'ha55ba566579b;
assign testcases[763] = 48'h434b97442a7c;
assign testcases[764] = 48'h21298842187c;
assign testcases[765] = 48'h11198811068b;
assign testcases[766] = 48'h00198811079b;
assign testcases[767] = 48'h00198810089b;
assign testcases[768] = 48'h00098800079b;
assign testcases[769] = 48'h00098800079b;
assign testcases[770] = 48'h00198800079b;
assign testcases[771] = 48'h00198800079b;
assign testcases[772] = 48'h00098800079b;
assign testcases[773] = 48'h00098800079b;
assign testcases[774] = 48'h332cc8421a9b;
assign testcases[775] = 48'h211ba821079b;
assign testcases[776] = 48'h110a9811079b;
assign testcases[777] = 48'h00098800079b;
assign testcases[778] = 48'h00098800079b;
assign testcases[779] = 48'h11198810079b;
assign testcases[780] = 48'h11198810179b;
assign testcases[781] = 48'h11098810079b;
assign testcases[782] = 48'h00098800079b;
assign testcases[783] = 48'h00098800079b;
assign testcases[784] = 48'h00098800079b;
assign testcases[785] = 48'h00099800079b;
assign testcases[786] = 48'h11177873199b;
assign testcases[787] = 48'h1008782106ab;
assign testcases[788] = 48'h10098800079b;
assign testcases[789] = 48'h221aa8741b6a;
assign testcases[790] = 48'h441988a6297a;
assign testcases[791] = 48'h661aa8d74a78;
assign testcases[792] = 48'h542bb8a63f43;
assign testcases[793] = 48'h212868733b77;
assign testcases[794] = 48'h11086811179b;
assign testcases[795] = 48'h11087811079b;
assign testcases[796] = 48'h11198811179b;
assign testcases[797] = 48'h11099811179b;
assign testcases[798] = 48'h121bf622179a;
assign testcases[799] = 48'h111ad711079b;
assign testcases[800] = 48'h111aa711079b;
assign testcases[801] = 48'h10099810079b;
assign testcases[802] = 48'h00098800079b;
assign testcases[803] = 48'h00098800079b;
assign testcases[804] = 48'h00098810079b;
assign testcases[805] = 48'h00098800079b;
assign testcases[806] = 48'h01099821189b;
assign testcases[807] = 48'h12198821189b;
assign testcases[808] = 48'h11198821079b;
assign testcases[809] = 48'h10099811079b;
assign testcases[810] = 48'h00099800079b;
assign testcases[811] = 48'h11184810179c;
assign testcases[812] = 48'h01097800079b;
assign testcases[813] = 48'h00098800079b;
assign testcases[814] = 48'h00199800079b;
assign testcases[815] = 48'h11199811079b;
assign testcases[816] = 48'h112a9811179b;
assign testcases[817] = 48'h11299811179a;
assign testcases[818] = 48'h01198811079b;
assign testcases[819] = 48'h00098811079b;
assign testcases[820] = 48'h00098800079b;
assign testcases[821] = 48'h00098800079b;
assign testcases[822] = 48'h02182910169c;
assign testcases[823] = 48'h01186800079b;
assign testcases[824] = 48'h01098800079b;
assign testcases[825] = 48'h00099800079b;
assign testcases[826] = 48'h01199811179b;
assign testcases[827] = 48'h0119981118aa;
assign testcases[828] = 48'h0009881117ab;
assign testcases[829] = 48'h00098801079b;
assign testcases[830] = 48'h11198811079b;
assign testcases[831] = 48'h11198811079b;
assign testcases[832] = 48'h00099800079b;
assign testcases[833] = 48'h00098800079b;
assign testcases[834] = 48'h11098801079b;
assign testcases[835] = 48'h11198811179c;
assign testcases[836] = 48'h11198711178b;
assign testcases[837] = 48'h875da3a697ab;
assign testcases[838] = 48'h977a85a6979b;
assign testcases[839] = 48'h987a87a6969b;
assign testcases[840] = 48'h987a98b7a79b;
assign testcases[841] = 48'ha77999b7989b;
assign testcases[842] = 48'h976889a787ab;
assign testcases[843] = 48'h977a8797979b;
assign testcases[844] = 48'h876a87a7969b;
assign testcases[845] = 48'h985999c7979b;
assign testcases[846] = 48'ha86898c7989b;
assign testcases[847] = 48'h975988b697ab;
assign testcases[848] = 48'h865a87a6979b;
assign testcases[849] = 48'h976a9796979c;
assign testcases[850] = 48'h873e83a6979c;
assign testcases[851] = 48'h875c95b6979b;
assign testcases[852] = 48'h865997b5989b;
assign testcases[853] = 48'h875989a5979b;
assign testcases[854] = 48'h865a7895979b;
assign testcases[855] = 48'h875a97a6979b;
assign testcases[856] = 48'h986998a6a79a;
assign testcases[857] = 48'h875889a6979b;
assign testcases[858] = 48'h876a88a697ab;
assign testcases[859] = 48'h875a87b6979b;
assign testcases[860] = 48'h875998b6969b;
assign testcases[861] = 48'h885898b6979b;
assign testcases[862] = 48'h986988b6979c;
assign testcases[863] = 48'h776a87c5d79c;
assign testcases[864] = 48'h776b85c5d69c;
assign testcases[865] = 48'h775b94c6c889;
assign testcases[866] = 48'h886998c7e89c;
assign testcases[867] = 48'h9a7987d6d7ac;
assign testcases[868] = 48'haa8988e6c79a;
assign testcases[869] = 48'hb8478cd7e7ac;
assign testcases[870] = 48'h99579bf5e78c;
assign testcases[871] = 48'h887a96e5e78b;
assign testcases[872] = 48'h886b94f6e69a;
assign testcases[873] = 48'h886997f6e7ab;
assign testcases[874] = 48'h887a96d5d99a;
assign testcases[875] = 48'ha89998d5d79d;
assign testcases[876] = 48'ha7578bc6e79c;
assign testcases[877] = 48'hb8bc94a676ca;
assign testcases[878] = 48'h887d9195779a;
assign testcases[879] = 48'ha9a7a8a6878b;
assign testcases[880] = 48'ha9889aa688ab;
assign testcases[881] = 48'h888b88a5889b;
assign testcases[882] = 48'h89797996868b;
assign testcases[883] = 48'h887b768576ab;
assign testcases[884] = 48'h877b8585779b;
assign testcases[885] = 48'h987d939686c9;
assign testcases[886] = 48'h997d9394979a;
assign testcases[887] = 48'haa9798a5878b;
assign testcases[888] = 48'ha9989aa5779a;
assign testcases[889] = 48'h899a8995779a;
assign testcases[890] = 48'h9a7999a5868c;
assign testcases[891] = 48'h898b86a597ad;
assign testcases[892] = 48'h698c84b497aa;
assign testcases[893] = 48'h798ba5a4889a;
assign testcases[894] = 48'hb9879aa6879c;
assign testcases[895] = 48'hc9889a96779b;
assign testcases[896] = 48'h88998995879a;
assign testcases[897] = 48'h897889b5968c;
assign testcases[898] = 48'h898b86b586ac;
assign testcases[899] = 48'h697c84a4879b;
assign testcases[900] = 48'h885c74c5d88d;
assign testcases[901] = 48'h885b74d6d69c;
assign testcases[902] = 48'h875b83e6c79a;
assign testcases[903] = 48'h977998e6d79c;
assign testcases[904] = 48'h997a87f7e69d;
assign testcases[905] = 48'h9a8998f7e899;
assign testcases[906] = 48'h88579be5f89b;
assign testcases[907] = 48'h113a882208ab;
assign testcases[908] = 48'h212a8712179b;
assign testcases[909] = 48'h111a8712179b;
assign testcases[910] = 48'h101a8801079b;
assign testcases[911] = 48'h00198801079b;
assign testcases[912] = 48'h00199801079b;
assign testcases[913] = 48'h00098800079b;
assign testcases[914] = 48'h00098800079b;
assign testcases[915] = 48'h00198800079b;
assign testcases[916] = 48'h00098800079b;
assign testcases[917] = 48'h00098800079b;
assign testcases[918] = 48'h00098800079b;
assign testcases[919] = 48'h11189811169b;
assign testcases[920] = 48'h00099800079b;
assign testcases[921] = 48'h00099800079b;
assign testcases[922] = 48'h00098800079b;
assign testcases[923] = 48'h00098800079b;
assign testcases[924] = 48'h00098800079b;
assign testcases[925] = 48'h00098800079b;
assign testcases[926] = 48'h00098800079b;
assign testcases[927] = 48'h00098800079b;
assign testcases[928] = 48'h00099800079b;
assign testcases[929] = 48'h11199811089b;
assign testcases[930] = 48'h100d771728c9;
assign testcases[931] = 48'h100c8802078b;
assign testcases[932] = 48'h100b8800079b;
assign testcases[933] = 48'h000a8800079b;
assign testcases[934] = 48'h00098800079b;
assign testcases[935] = 48'h00098800079b;
assign testcases[936] = 48'h00098800079b;
assign testcases[937] = 48'h00098800079b;
assign testcases[938] = 48'h00098800079b;
assign testcases[939] = 48'h00098800079b;
assign testcases[940] = 48'h00098800079b;
assign testcases[941] = 48'h00098800079b;
assign testcases[942] = 48'h3113772517e9;
assign testcases[943] = 48'h20068702179b;
assign testcases[944] = 48'h10088701079b;
assign testcases[945] = 48'h00099800079b;
assign testcases[946] = 48'h000a9800079b;
assign testcases[947] = 48'h000a8800079b;
assign testcases[948] = 48'h00098800079b;
assign testcases[949] = 48'h00098800079b;
assign testcases[950] = 48'h00098800079b;
assign testcases[951] = 48'h00098800079b;
assign testcases[952] = 48'h00098800079b;
assign testcases[953] = 48'h00098800079b;
assign testcases[954] = 48'h441e8822369f;
assign testcases[955] = 48'h110b9800179b;
assign testcases[956] = 48'h10099800079b;
assign testcases[957] = 48'h00098800079b;
assign testcases[958] = 48'h00098800079b;
assign testcases[959] = 48'h00098800079b;
assign testcases[960] = 48'h00098800079b;
assign testcases[961] = 48'h00098800079b;
assign testcases[962] = 48'h00098800079b;
assign testcases[963] = 48'h00098800079b;
assign testcases[964] = 48'h00098800079b;
assign testcases[965] = 48'h00098800079b;
assign testcases[966] = 48'h00098800079b;
assign testcases[967] = 48'h00099800079b;
assign testcases[968] = 48'h00098800079b;
assign testcases[969] = 48'h226cf8974008;
assign testcases[970] = 48'h114bc822178c;
assign testcases[971] = 48'h111aa710079b;
assign testcases[972] = 48'h001a9710079b;
assign testcases[973] = 48'h00098700079b;
assign testcases[974] = 48'h0009880107ab;
assign testcases[975] = 48'h00098801079b;
assign testcases[976] = 48'h00098801078b;
assign testcases[977] = 48'h00098800079b;
assign testcases[978] = 48'h00098800079b;
assign testcases[979] = 48'h00098800079b;
assign testcases[980] = 48'h00098800079b;
assign testcases[981] = 48'h00098800079b;
assign testcases[982] = 48'h00098800079b;
assign testcases[983] = 48'h00098800079b;
assign testcases[984] = 48'h00198811079b;
assign testcases[985] = 48'h97797a69879a;
assign testcases[986] = 48'ha769887998ac;
assign testcases[987] = 48'ha7798869a79c;
assign testcases[988] = 48'ha88a8879979a;
assign testcases[989] = 48'ha87a977986ab;
assign testcases[990] = 48'hb8699779878c;
assign testcases[991] = 48'ha8789879878b;
assign testcases[992] = 48'h9879977987aa;
assign testcases[993] = 48'ha8698879989c;
assign testcases[994] = 48'ha8799878979c;
assign testcases[995] = 48'ha87a8868979a;
assign testcases[996] = 48'h977a8869779b;
assign testcases[997] = 48'h9779886a77ac;
assign testcases[998] = 48'h9768877a778c;
assign testcases[999] = 48'h977a7a68789a;


  
  localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
  wire [$clog2(CLASS_CNT)-1:0] prediction;

  // Instantiate module under test
 Har_tnn1_tnnseq #(
 ) dut (
    .data(data),
    .clk(clk),
    .rst(rst),
    .prediction(prediction)
  );
  
  always #halfT clk <= ~clk;

  integer i,j;
  initial begin
    for(i=0;i<TEST_CNT;i=i+1)
        runtestcase(i);
    $finish;
  end

  task runtestcase(input integer i); begin
    data <= testcases[i];
    rst <= 1;
    clk <= 0;
    #period
    rst <= 0;
    #period
    #((FEAT_CNT+HIDDEN_CNT-1)*period)
    for (j = 0; j < CLASS_CNT; j=j+1) begin
        $write("%d ,",dut.tnn.scores[j*7+:7]);
    end
    $display("");
    /* $display("%h",dut.tnn.scores); */
  end
  endtask

endmodule
