













module cardio_bnn1_bnnroperm #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 760'b1110000110110101010011010111011011101101110101001000010100111010010000101110111100001011001111001101101101101110100010000000110011110010111001001010101011001011110001100011100000111011101100100010110110011000111100101110101000101000001001000110000011000001100011000101101000000110000000001100100011000101100001110001000010110001010011010101010010010100000010100100111000100000010000001110101111010110010101001001010001000111101011000101100010010010110100011010010000100011101000001101111110010010100111111100100011000000111101110100001011000010110101111110110100011010011101000000010000001100000001010010000111100100000100101010000000001101110100101010101011100111000111111000001110100111001010111001010011101101011010101100110010001111011000111101000110101011 ;
  localparam Weights1 = 120'b100111001101000001001001110101000100000111111001000100000010111111100110010111111111110100010000001010101000111001011111 ;

  romesh_seq #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
