












module winequality_white_bnn_seq #(

parameter N = 11,
parameter M = 40,
parameter B = 4,
parameter C = 7,
parameter Ts = 5


  ) (
  input clk,
  input rst,
  input [N*B-1:0] data,
  output [$clog2(C)-1:0] klass
  );

  localparam Weights0 = 440'b01011011001001010110011000111111100001101110011110111101111010000011000010100110111100010000110010110011100101010111010001001000111000101011010101001110010111011110101100111011111000110011011010110110011111001000001111001101001001101000010110100001111111101110001001001000111100001010010111011000101010001111011111100101110010110001011100100001001001110010100011000000000001001011010100011010101110001001110001001010111111100000111001011000 ;
  localparam Weights1 = 280'b0110101101111010110110010101001100000000111001110111011111111000110100011011000011101011011100101111000011010111101100001100101101000010001100000101011110110000111010110111001011111000110101111101100011101011011100101111110011000111101100011110001101010011010011001100000001110011 ;

  localparam SumL = $clog2(M+1);
  wire [SumL*C-1:0] sums;

  seqlego #(.N(N),.B(B),.M(M),.C(C),.Weights0(Weights0),.Weights1(Weights1)) layers (
    .clk(clk),
    .rst(rst),
    .data(data),
    .out(sums)
  );

  argmax #(.N(C),.I($clog2(C)),.K(SumL)) result (
     .inx(sums),
     .outimax(klass)
  );

endmodule
