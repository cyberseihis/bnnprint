`timescale 1us/1ns









module tbwinequality_white_bs #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1000


)();

  
  reg [FEAT_BITS*FEAT_CNT-1:0] sample;
  wire [FEAT_BITS*FEAT_CNT-1:0] testcases [TEST_CNT-1:0];
  reg rst;
  reg clk;
  parameter Nsperiod=50000;
  localparam period=Nsperiod/500;
  localparam halfPeriod=period/2;


assign testcases[0] = 44'h53352264442;
assign testcases[1] = 44'h43302152854;
assign testcases[2] = 44'h73422232845;
assign testcases[3] = 44'h52322373735;
assign testcases[4] = 44'h52322373735;
assign testcases[5] = 44'h73422232845;
assign testcases[6] = 44'h44222252754;
assign testcases[7] = 44'h53352264442;
assign testcases[8] = 44'h43302152854;
assign testcases[9] = 44'h72402142748;
assign testcases[10] = 44'h7340112146a;
assign testcases[11] = 44'h72411142664;
assign testcases[12] = 44'h62401122787;
assign testcases[13] = 44'h41402351c6b;
assign testcases[14] = 44'h75651264484;
assign testcases[15] = 44'h41401141869;
assign testcases[16] = 44'h46002232834;
assign testcases[17] = 44'h4950122193c;
assign testcases[18] = 44'h64401161669;
assign testcases[19] = 44'h44122253754;
assign testcases[20] = 44'h4950122193c;
assign testcases[21] = 44'h44411131728;
assign testcases[22] = 44'h53402242b56;
assign testcases[23] = 44'h69103162553;
assign testcases[24] = 44'h43402152a55;
assign testcases[25] = 44'h53322393856;
assign testcases[26] = 44'h53302252b45;
assign testcases[27] = 44'h53422253a66;
assign testcases[28] = 44'h63502151759;
assign testcases[29] = 44'h5430124169b;
assign testcases[30] = 44'h73422153765;
assign testcases[31] = 44'h71302012b36;
assign testcases[32] = 44'h63302232747;
assign testcases[33] = 44'h41302242a53;
assign testcases[34] = 44'h33242163936;
assign testcases[35] = 44'h5340314174c;
assign testcases[36] = 44'h45212152825;
assign testcases[37] = 44'h54302251618;
assign testcases[38] = 44'h53442254732;
assign testcases[39] = 44'h53442254732;
assign testcases[40] = 44'h42408362634;
assign testcases[41] = 44'h43418352624;
assign testcases[42] = 44'h54323163645;
assign testcases[43] = 44'h43302252764;
assign testcases[44] = 44'h42302252864;
assign testcases[45] = 44'h62302262665;
assign testcases[46] = 44'h46313372865;
assign testcases[47] = 44'h46213372865;
assign testcases[48] = 44'h54323163645;
assign testcases[49] = 44'h52313252955;
assign testcases[50] = 44'h5230326194a;
assign testcases[51] = 44'h43303241978;
assign testcases[52] = 44'h41302131947;
assign testcases[53] = 44'h42302241927;
assign testcases[54] = 44'h52607252533;
assign testcases[55] = 44'h53301271668;
assign testcases[56] = 44'h52332283554;
assign testcases[57] = 44'h32332353832;
assign testcases[58] = 44'h45112132636;
assign testcases[59] = 44'h62301242925;
assign testcases[60] = 44'h52214242542;
assign testcases[61] = 44'h32332353832;
assign testcases[62] = 44'h56101151426;
assign testcases[63] = 44'h45112132636;
assign testcases[64] = 44'h53301242646;
assign testcases[65] = 44'h44003242763;
assign testcases[66] = 44'h4321114175c;
assign testcases[67] = 44'h43102462645;
assign testcases[68] = 44'h42302232987;
assign testcases[69] = 44'h63322143624;
assign testcases[70] = 44'h43422393653;
assign testcases[71] = 44'h53212393974;
assign testcases[72] = 44'h33313273e95;
assign testcases[73] = 44'h72402022353;
assign testcases[74] = 44'h42302232987;
assign testcases[75] = 44'h63322143624;
assign testcases[76] = 44'h5230223183c;
assign testcases[77] = 44'h5430212198a;
assign testcases[78] = 44'h62323133363;
assign testcases[79] = 44'h47312142833;
assign testcases[80] = 44'h52302242aa7;
assign testcases[81] = 44'h52342364773;
assign testcases[82] = 44'h54213362745;
assign testcases[83] = 44'h52322273944;
assign testcases[84] = 44'h55632353642;
assign testcases[85] = 44'h56632353642;
assign testcases[86] = 44'h55632353542;
assign testcases[87] = 44'h53332473754;
assign testcases[88] = 44'h55632353642;
assign testcases[89] = 44'h56632353642;
assign testcases[90] = 44'h55632353542;
assign testcases[91] = 44'h43422493653;
assign testcases[92] = 44'h5330135183c;
assign testcases[93] = 44'h5230135184c;
assign testcases[94] = 44'h61301351749;
assign testcases[95] = 44'h53332393543;
assign testcases[96] = 44'h34642163652;
assign testcases[97] = 44'h73301131339;
assign testcases[98] = 44'h94421033215;
assign testcases[99] = 44'h34642163652;
assign testcases[100] = 44'h63432373443;
assign testcases[101] = 44'h51322363a44;
assign testcases[102] = 44'h32232363934;
assign testcases[103] = 44'h64442264443;
assign testcases[104] = 44'h63432373443;
assign testcases[105] = 44'h51332243723;
assign testcases[106] = 44'h51322363a44;
assign testcases[107] = 44'h52341364673;
assign testcases[108] = 44'h52341364673;
assign testcases[109] = 44'h54302272876;
assign testcases[110] = 44'h41523363232;
assign testcases[111] = 44'h53442294562;
assign testcases[112] = 44'h54532473453;
assign testcases[113] = 44'h45322253753;
assign testcases[114] = 44'h45322253753;
assign testcases[115] = 44'h36003032d34;
assign testcases[116] = 44'h34212151949;
assign testcases[117] = 44'h5140113174a;
assign testcases[118] = 44'h54532473453;
assign testcases[119] = 44'h54532373553;
assign testcases[120] = 44'h34012132756;
assign testcases[121] = 44'h63332253462;
assign testcases[122] = 44'h61322252824;
assign testcases[123] = 44'h52312152833;
assign testcases[124] = 44'h41504262735;
assign testcases[125] = 44'h42301351858;
assign testcases[126] = 44'h65221242646;
assign testcases[127] = 44'h43321373b64;
assign testcases[128] = 44'h43512362877;
assign testcases[129] = 44'h43512262977;
assign testcases[130] = 44'h33221022a37;
assign testcases[131] = 44'h43321373b64;
assign testcases[132] = 44'h45431393773;
assign testcases[133] = 44'h43341273853;
assign testcases[134] = 44'h53221373762;
assign testcases[135] = 44'h43341263864;
assign testcases[136] = 44'h72401242637;
assign testcases[137] = 44'h55622353642;
assign testcases[138] = 44'h52301231667;
assign testcases[139] = 44'h7340113276a;
assign testcases[140] = 44'h44302132846;
assign testcases[141] = 44'h55622353642;
assign testcases[142] = 44'h62401242767;
assign testcases[143] = 44'h72411132764;
assign testcases[144] = 44'h72401132668;
assign testcases[145] = 44'h43401241437;
assign testcases[146] = 44'h31302361835;
assign testcases[147] = 44'h48112132a33;
assign testcases[148] = 44'h44311131a7a;
assign testcases[149] = 44'h53312142434;
assign testcases[150] = 44'h62422252629;
assign testcases[151] = 44'h62422353645;
assign testcases[152] = 44'h53312142434;
assign testcases[153] = 44'h52402231646;
assign testcases[154] = 44'h724221235c4;
assign testcases[155] = 44'h63433373242;
assign testcases[156] = 44'h63433373242;
assign testcases[157] = 44'h4420124184b;
assign testcases[158] = 44'h2600124192b;
assign testcases[159] = 44'h2600124192b;
assign testcases[160] = 44'h4420124184b;
assign testcases[161] = 44'h42532163433;
assign testcases[162] = 44'h44312132837;
assign testcases[163] = 44'h63433373242;
assign testcases[164] = 44'h43332373654;
assign testcases[165] = 44'h52332463655;
assign testcases[166] = 44'h73422273674;
assign testcases[167] = 44'h4620113154c;
assign testcases[168] = 44'h63322153563;
assign testcases[169] = 44'h95521043215;
assign testcases[170] = 44'h5340325166c;
assign testcases[171] = 44'h62402131638;
assign testcases[172] = 44'h66401031539;
assign testcases[173] = 44'h42411241929;
assign testcases[174] = 44'h63342264586;
assign testcases[175] = 44'h52421352619;
assign testcases[176] = 44'h5451212154c;
assign testcases[177] = 44'h32332363834;
assign testcases[178] = 44'h39102042622;
assign testcases[179] = 44'h43312262793;
assign testcases[180] = 44'h44312262783;
assign testcases[181] = 44'h54102362543;
assign testcases[182] = 44'h53452364352;
assign testcases[183] = 44'h53432383774;
assign testcases[184] = 44'h53532383483;
assign testcases[185] = 44'h53532483483;
assign testcases[186] = 44'h43421363675;
assign testcases[187] = 44'h33211242658;
assign testcases[188] = 44'h5731114187c;
assign testcases[189] = 44'h43322373562;
assign testcases[190] = 44'h43322373562;
assign testcases[191] = 44'h53452364352;
assign testcases[192] = 44'h53322142439;
assign testcases[193] = 44'h41312242944;
assign testcases[194] = 44'h43419462443;
assign testcases[195] = 44'h43419462433;
assign testcases[196] = 44'h43419462433;
assign testcases[197] = 44'h53222383652;
assign testcases[198] = 44'h54232373652;
assign testcases[199] = 44'h53222383652;
assign testcases[200] = 44'h53342373653;
assign testcases[201] = 44'h54232373652;
assign testcases[202] = 44'h57332383754;
assign testcases[203] = 44'h5333125296a;
assign testcases[204] = 44'h33302242856;
assign testcases[205] = 44'h42532253642;
assign testcases[206] = 44'h51322243723;
assign testcases[207] = 44'ha6812143455;
assign testcases[208] = 44'h583011329a6;
assign testcases[209] = 44'h453021627a4;
assign testcases[210] = 44'h33221122926;
assign testcases[211] = 44'h52401241978;
assign testcases[212] = 44'h51322243723;
assign testcases[213] = 44'h41312242a34;
assign testcases[214] = 44'h43201241848;
assign testcases[215] = 44'h33222353934;
assign testcases[216] = 44'h63321262528;
assign testcases[217] = 44'h33222353934;
assign testcases[218] = 44'h33242364944;
assign testcases[219] = 44'h62321262528;
assign testcases[220] = 44'h63321262528;
assign testcases[221] = 44'h59223263463;
assign testcases[222] = 44'h43201241848;
assign testcases[223] = 44'h42302252a33;
assign testcases[224] = 44'h47202252a66;
assign testcases[225] = 44'h53442254932;
assign testcases[226] = 44'h41302272b54;
assign testcases[227] = 44'h533224a3763;
assign testcases[228] = 44'h41302272b54;
assign testcases[229] = 44'h53442254932;
assign testcases[230] = 44'h59123153942;
assign testcases[231] = 44'h73422273954;
assign testcases[232] = 44'h73421373954;
assign testcases[233] = 44'h52432373543;
assign testcases[234] = 44'h52432373543;
assign testcases[235] = 44'h52432373543;
assign testcases[236] = 44'h52432373543;
assign testcases[237] = 44'h57332383854;
assign testcases[238] = 44'h53601241948;
assign testcases[239] = 44'h43241163b84;
assign testcases[240] = 44'h54232374742;
assign testcases[241] = 44'h64321132656;
assign testcases[242] = 44'h52401131639;
assign testcases[243] = 44'h53312382874;
assign testcases[244] = 44'h55532253642;
assign testcases[245] = 44'h423011929b9;
assign testcases[246] = 44'h5230115167c;
assign testcases[247] = 44'h32301131837;
assign testcases[248] = 44'h32301121837;
assign testcases[249] = 44'h45121143a45;
assign testcases[250] = 44'h32312273f95;
assign testcases[251] = 44'h73243273455;
assign testcases[252] = 44'h55532253642;
assign testcases[253] = 44'h33411041c4a;
assign testcases[254] = 44'h33402262763;
assign testcases[255] = 44'h43401252974;
assign testcases[256] = 44'h44311032848;
assign testcases[257] = 44'h44311032848;
assign testcases[258] = 44'h4240114195a;
assign testcases[259] = 44'h34401021829;
assign testcases[260] = 44'h51312242946;
assign testcases[261] = 44'h53452254352;
assign testcases[262] = 44'h53421132726;
assign testcases[263] = 44'h53432483574;
assign testcases[264] = 44'h43301161657;
assign testcases[265] = 44'h53452254352;
assign testcases[266] = 44'h54322263853;
assign testcases[267] = 44'h28122252974;
assign testcases[268] = 44'h28122252974;
assign testcases[269] = 44'h28122252974;
assign testcases[270] = 44'h54322263853;
assign testcases[271] = 44'h28122252974;
assign testcases[272] = 44'h33332253833;
assign testcases[273] = 44'h48312242833;
assign testcases[274] = 44'h53522383574;
assign testcases[275] = 44'h42422363675;
assign testcases[276] = 44'h42422363675;
assign testcases[277] = 44'h63402021257;
assign testcases[278] = 44'h54302121557;
assign testcases[279] = 44'h5351114189b;
assign testcases[280] = 44'h5331114173c;
assign testcases[281] = 44'h4461124187b;
assign testcases[282] = 44'h56412272586;
assign testcases[283] = 44'h44342373753;
assign testcases[284] = 44'h54242274652;
assign testcases[285] = 44'h54222363552;
assign testcases[286] = 44'h43342373754;
assign testcases[287] = 44'h52432373453;
assign testcases[288] = 44'h52432373453;
assign testcases[289] = 44'h52432373453;
assign testcases[290] = 44'h52432373453;
assign testcases[291] = 44'h31312352c46;
assign testcases[292] = 44'h63453374343;
assign testcases[293] = 44'h43222153a85;
assign testcases[294] = 44'h88403263731;
assign testcases[295] = 44'h44302262964;
assign testcases[296] = 44'h75722263574;
assign testcases[297] = 44'h52412472778;
assign testcases[298] = 44'h61432453745;
assign testcases[299] = 44'h41502142646;
assign testcases[300] = 44'h45003231887;
assign testcases[301] = 44'h72302122636;
assign testcases[302] = 44'h45003231887;
assign testcases[303] = 44'h33202261948;
assign testcases[304] = 44'h55222262745;
assign testcases[305] = 44'h55222262745;
assign testcases[306] = 44'h55212262745;
assign testcases[307] = 44'h55212262745;
assign testcases[308] = 44'h44311252746;
assign testcases[309] = 44'h44311252746;
assign testcases[310] = 44'h44301131a99;
assign testcases[311] = 44'h27121261c5c;
assign testcases[312] = 44'h63412253945;
assign testcases[313] = 44'h34211362885;
assign testcases[314] = 44'h34211362875;
assign testcases[315] = 44'h53606242543;
assign testcases[316] = 44'h53311252737;
assign testcases[317] = 44'h43321252736;
assign testcases[318] = 44'h33521152c49;
assign testcases[319] = 44'h41211022c75;
assign testcases[320] = 44'h30202122d76;
assign testcases[321] = 44'h43321252736;
assign testcases[322] = 44'h53311252737;
assign testcases[323] = 44'h53421252636;
assign testcases[324] = 44'h75502172469;
assign testcases[325] = 44'h633127b2776;
assign testcases[326] = 44'h63441283375;
assign testcases[327] = 44'h44211252785;
assign testcases[328] = 44'h43342373754;
assign testcases[329] = 44'h52401232756;
assign testcases[330] = 44'h4431123197c;
assign testcases[331] = 44'h53311252737;
assign testcases[332] = 44'h4230113183a;
assign testcases[333] = 44'h43321253645;
assign testcases[334] = 44'h33311132837;
assign testcases[335] = 44'h4230113183a;
assign testcases[336] = 44'h42301141948;
assign testcases[337] = 44'h33332363843;
assign testcases[338] = 44'h33402152b66;
assign testcases[339] = 44'h42302352ac6;
assign testcases[340] = 44'h62422153763;
assign testcases[341] = 44'h63302142765;
assign testcases[342] = 44'h43422253753;
assign testcases[343] = 44'h245122528a5;
assign testcases[344] = 44'h235123528a5;
assign testcases[345] = 44'h51312252834;
assign testcases[346] = 44'h34101121958;
assign testcases[347] = 44'h42442454742;
assign testcases[348] = 44'h62432243655;
assign testcases[349] = 44'h61432353655;
assign testcases[350] = 44'h413023518a9;
assign testcases[351] = 44'h5442125251a;
assign testcases[352] = 44'h34303142654;
assign testcases[353] = 44'h5442125251a;
assign testcases[354] = 44'h35412292874;
assign testcases[355] = 44'h52433373233;
assign testcases[356] = 44'h52433373233;
assign testcases[357] = 44'h443021626a4;
assign testcases[358] = 44'ha2402152446;
assign testcases[359] = 44'h53311262777;
assign testcases[360] = 44'h43342363856;
assign testcases[361] = 44'h54102132642;
assign testcases[362] = 44'h51312242a34;
assign testcases[363] = 44'h52433373233;
assign testcases[364] = 44'h51401132b49;
assign testcases[365] = 44'h33311241a9b;
assign testcases[366] = 44'h32304252b77;
assign testcases[367] = 44'h54202252644;
assign testcases[368] = 44'h63502262787;
assign testcases[369] = 44'h55332122719;
assign testcases[370] = 44'h54202252644;
assign testcases[371] = 44'h63502262787;
assign testcases[372] = 44'h4d202172965;
assign testcases[373] = 44'h53302252653;
assign testcases[374] = 44'h24201131b3c;
assign testcases[375] = 44'h24201131b3c;
assign testcases[376] = 44'h44301141956;
assign testcases[377] = 44'h52402132645;
assign testcases[378] = 44'h34502152785;
assign testcases[379] = 44'h44301141956;
assign testcases[380] = 44'h52402132645;
assign testcases[381] = 44'h53332363663;
assign testcases[382] = 44'h64322153663;
assign testcases[383] = 44'h53302252653;
assign testcases[384] = 44'h34411141a39;
assign testcases[385] = 44'h24201131b3c;
assign testcases[386] = 44'h21501141b37;
assign testcases[387] = 44'h45311492685;
assign testcases[388] = 44'h42312252a44;
assign testcases[389] = 44'h53441363773;
assign testcases[390] = 44'h53441363773;
assign testcases[391] = 44'h44301121647;
assign testcases[392] = 44'h47121143956;
assign testcases[393] = 44'h5340112156b;
assign testcases[394] = 44'h55532363742;
assign testcases[395] = 44'h53101562745;
assign testcases[396] = 44'h73401231539;
assign testcases[397] = 44'h42401241b59;
assign testcases[398] = 44'h33342364944;
assign testcases[399] = 44'h4241123184a;
assign testcases[400] = 44'h42401241b59;
assign testcases[401] = 44'h55532363742;
assign testcases[402] = 44'h44103142763;
assign testcases[403] = 44'h53342394562;
assign testcases[404] = 44'h5231126188c;
assign testcases[405] = 44'h53101562745;
assign testcases[406] = 44'h33311231a3c;
assign testcases[407] = 44'h56202142754;
assign testcases[408] = 44'h41402142866;
assign testcases[409] = 44'h73401231539;
assign testcases[410] = 44'h53451254453;
assign testcases[411] = 44'h533312538b4;
assign testcases[412] = 44'h52401231656;
assign testcases[413] = 44'h52401231656;
assign testcases[414] = 44'h53451254453;
assign testcases[415] = 44'h533312538b4;
assign testcases[416] = 44'h62302132725;
assign testcases[417] = 44'h53222373653;
assign testcases[418] = 44'h62302132725;
assign testcases[419] = 44'h64302252966;
assign testcases[420] = 44'h5231125163c;
assign testcases[421] = 44'h52322283866;
assign testcases[422] = 44'h52322283866;
assign testcases[423] = 44'h52322283866;
assign testcases[424] = 44'h52422363966;
assign testcases[425] = 44'h52322283866;
assign testcases[426] = 44'h52322283866;
assign testcases[427] = 44'h53532373544;
assign testcases[428] = 44'h62302132543;
assign testcases[429] = 44'h54532373653;
assign testcases[430] = 44'h53532373544;
assign testcases[431] = 44'h44102132735;
assign testcases[432] = 44'h61302482775;
assign testcases[433] = 44'h57105152573;
assign testcases[434] = 44'h5232124295b;
assign testcases[435] = 44'h52411132a5b;
assign testcases[436] = 44'h43302182875;
assign testcases[437] = 44'h4130137198b;
assign testcases[438] = 44'h61302482775;
assign testcases[439] = 44'h44002142863;
assign testcases[440] = 44'h42401131879;
assign testcases[441] = 44'h45211152896;
assign testcases[442] = 44'h33301341a8d;
assign testcases[443] = 44'h47432393863;
assign testcases[444] = 44'h53351253728;
assign testcases[445] = 44'h54331122839;
assign testcases[446] = 44'h33302251c4b;
assign testcases[447] = 44'h45232143a65;
assign testcases[448] = 44'h45232143a65;
assign testcases[449] = 44'h43302242b66;
assign testcases[450] = 44'h58223163563;
assign testcases[451] = 44'h42201242845;
assign testcases[452] = 44'h36112162b57;
assign testcases[453] = 44'h33302242a56;
assign testcases[454] = 44'h43302242b66;
assign testcases[455] = 44'h45232143a65;
assign testcases[456] = 44'h4230113183d;
assign testcases[457] = 44'h52322143364;
assign testcases[458] = 44'h35302282895;
assign testcases[459] = 44'h45322593951;
assign testcases[460] = 44'h52322143364;
assign testcases[461] = 44'h53342263743;
assign testcases[462] = 44'h33232363934;
assign testcases[463] = 44'h54202122734;
assign testcases[464] = 44'h55632463652;
assign testcases[465] = 44'h42623243342;
assign testcases[466] = 44'h51321353744;
assign testcases[467] = 44'h54202122734;
assign testcases[468] = 44'h55632463652;
assign testcases[469] = 44'h53542364564;
assign testcases[470] = 44'h75731163493;
assign testcases[471] = 44'h453112726a5;
assign testcases[472] = 44'h4330113184c;
assign testcases[473] = 44'h51311252954;
assign testcases[474] = 44'h31211232834;
assign testcases[475] = 44'h53531383574;
assign testcases[476] = 44'h6330124143b;
assign testcases[477] = 44'h52301242666;
assign testcases[478] = 44'h57103162473;
assign testcases[479] = 44'h42302462966;
assign testcases[480] = 44'h46322263773;
assign testcases[481] = 44'h34402241957;
assign testcases[482] = 44'h33232253944;
assign testcases[483] = 44'h46322263773;
assign testcases[484] = 44'h4531f473874;
assign testcases[485] = 44'h42401242b64;
assign testcases[486] = 44'h31401242b54;
assign testcases[487] = 44'h44301231647;
assign testcases[488] = 44'h63302362996;
assign testcases[489] = 44'h63322363642;
assign testcases[490] = 44'h5330102154b;
assign testcases[491] = 44'h5240112183c;
assign testcases[492] = 44'h62321263745;
assign testcases[493] = 44'h42301161789;
assign testcases[494] = 44'h52411132977;
assign testcases[495] = 44'h3612116195c;
assign testcases[496] = 44'h55632473552;
assign testcases[497] = 44'h5230125186c;
assign testcases[498] = 44'h34301162885;
assign testcases[499] = 44'h55632473552;
assign testcases[500] = 44'h53542374554;
assign testcases[501] = 44'h52631363654;
assign testcases[502] = 44'h43301072775;
assign testcases[503] = 44'h43301072775;
assign testcases[504] = 44'h62332253562;
assign testcases[505] = 44'h62332253562;
assign testcases[506] = 44'h57314052462;
assign testcases[507] = 44'h33302262d65;
assign testcases[508] = 44'h38311351a4a;
assign testcases[509] = 44'h33302262d65;
assign testcases[510] = 44'h43102352745;
assign testcases[511] = 44'h6430206164b;
assign testcases[512] = 44'h53311252678;
assign testcases[513] = 44'h64301121728;
assign testcases[514] = 44'h63321242736;
assign testcases[515] = 44'h44302162956;
assign testcases[516] = 44'h52402352543;
assign testcases[517] = 44'h61402352476;
assign testcases[518] = 44'h31302131a87;
assign testcases[519] = 44'h5433201273a;
assign testcases[520] = 44'h623010525a5;
assign testcases[521] = 44'h623010525a5;
assign testcases[522] = 44'h53401131539;
assign testcases[523] = 44'h34301131538;
assign testcases[524] = 44'h34401021929;
assign testcases[525] = 44'h34415152543;
assign testcases[526] = 44'h5441101156c;
assign testcases[527] = 44'h4320124194c;
assign testcases[528] = 44'h24001141a2b;
assign testcases[529] = 44'h32511142c48;
assign testcases[530] = 44'h40312232ab4;
assign testcases[531] = 44'h42518352533;
assign testcases[532] = 44'h63333363453;
assign testcases[533] = 44'h63333363453;
assign testcases[534] = 44'h63333363453;
assign testcases[535] = 44'h64542364553;
assign testcases[536] = 44'h64542364553;
assign testcases[537] = 44'h63333363453;
assign testcases[538] = 44'h43302122966;
assign testcases[539] = 44'h53212273984;
assign testcases[540] = 44'h44321063b69;
assign testcases[541] = 44'h56622473642;
assign testcases[542] = 44'h34302162995;
assign testcases[543] = 44'h43421252775;
assign testcases[544] = 44'h53232363753;
assign testcases[545] = 44'h41201252b75;
assign testcases[546] = 44'h43221263b84;
assign testcases[547] = 44'h6240203285a;
assign testcases[548] = 44'h42302242b56;
assign testcases[549] = 44'h56622473642;
assign testcases[550] = 44'h53532263564;
assign testcases[551] = 44'h83301231339;
assign testcases[552] = 44'h6330124143b;
assign testcases[553] = 44'h53532263564;
assign testcases[554] = 44'h6330124143b;
assign testcases[555] = 44'h83301231339;
assign testcases[556] = 44'h74732163484;
assign testcases[557] = 44'h45202152956;
assign testcases[558] = 44'h32232363834;
assign testcases[559] = 44'h544123514ab;
assign testcases[560] = 44'h424222536a5;
assign testcases[561] = 44'h35102242855;
assign testcases[562] = 44'h64323263583;
assign testcases[563] = 44'h632021525a6;
assign testcases[564] = 44'h57313262743;
assign testcases[565] = 44'h62422133655;
assign testcases[566] = 44'h54332012639;
assign testcases[567] = 44'h33502352575;
assign testcases[568] = 44'h43502352575;
assign testcases[569] = 44'h43311262794;
assign testcases[570] = 44'h65632473542;
assign testcases[571] = 44'h43311141949;
assign testcases[572] = 44'h44542264562;
assign testcases[573] = 44'h5231135163c;
assign testcases[574] = 44'h6230125174a;
assign testcases[575] = 44'h72302372656;
assign testcases[576] = 44'h72302372656;
assign testcases[577] = 44'h5231135163c;
assign testcases[578] = 44'h43311141949;
assign testcases[579] = 44'h35311251a3b;
assign testcases[580] = 44'h65632473542;
assign testcases[581] = 44'h32212142934;
assign testcases[582] = 44'h53212262625;
assign testcases[583] = 44'h63222133234;
assign testcases[584] = 44'h43302252a55;
assign testcases[585] = 44'h63222133234;
assign testcases[586] = 44'h63322253652;
assign testcases[587] = 44'h44201252b57;
assign testcases[588] = 44'h53301242a57;
assign testcases[589] = 44'h52311152774;
assign testcases[590] = 44'h54532053343;
assign testcases[591] = 44'h52401342957;
assign testcases[592] = 44'h55322153764;
assign testcases[593] = 44'h46101051417;
assign testcases[594] = 44'h46101051417;
assign testcases[595] = 44'h43402052b56;
assign testcases[596] = 44'h55322153764;
assign testcases[597] = 44'h53411142747;
assign testcases[598] = 44'h33331242956;
assign testcases[599] = 44'h52401121599;
assign testcases[600] = 44'h43308262664;
assign testcases[601] = 44'h53402241237;
assign testcases[602] = 44'h46101051417;
assign testcases[603] = 44'h46101051417;
assign testcases[604] = 44'h43502252475;
assign testcases[605] = 44'h43502252475;
assign testcases[606] = 44'h53322263a34;
assign testcases[607] = 44'h53322263a34;
assign testcases[608] = 44'h43242364954;
assign testcases[609] = 44'h65312133b97;
assign testcases[610] = 44'h4431124188b;
assign testcases[611] = 44'h63411032538;
assign testcases[612] = 44'h62732253432;
assign testcases[613] = 44'h62732253432;
assign testcases[614] = 44'h62732253432;
assign testcases[615] = 44'h62732253432;
assign testcases[616] = 44'h6430113178a;
assign testcases[617] = 44'h63302372757;
assign testcases[618] = 44'h63302372757;
assign testcases[619] = 44'h62302252654;
assign testcases[620] = 44'h46444384773;
assign testcases[621] = 44'h43424363253;
assign testcases[622] = 44'h24112152976;
assign testcases[623] = 44'h53302021759;
assign testcases[624] = 44'h34103142863;
assign testcases[625] = 44'h43331342948;
assign testcases[626] = 44'h68124163943;
assign testcases[627] = 44'h54212283774;
assign testcases[628] = 44'h54212283774;
assign testcases[629] = 44'h34301131776;
assign testcases[630] = 44'h52442254742;
assign testcases[631] = 44'h52442254742;
assign testcases[632] = 44'h53311152887;
assign testcases[633] = 44'h33232273944;
assign testcases[634] = 44'h41311252a57;
assign testcases[635] = 44'h31211252b57;
assign testcases[636] = 44'h41311252a47;
assign testcases[637] = 44'h63232153673;
assign testcases[638] = 44'h34112372896;
assign testcases[639] = 44'h34112372896;
assign testcases[640] = 44'h32302241958;
assign testcases[641] = 44'h43232273843;
assign testcases[642] = 44'h42332463956;
assign testcases[643] = 44'h43332263944;
assign testcases[644] = 44'h43332263944;
assign testcases[645] = 44'h43222263843;
assign testcases[646] = 44'h44702052574;
assign testcases[647] = 44'h60332353633;
assign testcases[648] = 44'h34112272695;
assign testcases[649] = 44'h53333274563;
assign testcases[650] = 44'h53333274563;
assign testcases[651] = 44'h53333274563;
assign testcases[652] = 44'h53333274563;
assign testcases[653] = 44'h33332253944;
assign testcases[654] = 44'h424024519a9;
assign testcases[655] = 44'h6331124264b;
assign testcases[656] = 44'h83311132539;
assign testcases[657] = 44'h54212152846;
assign testcases[658] = 44'h43212271839;
assign testcases[659] = 44'h53201782655;
assign testcases[660] = 44'h53302132634;
assign testcases[661] = 44'h5333135295b;
assign testcases[662] = 44'h58124173a53;
assign testcases[663] = 44'h53302132634;
assign testcases[664] = 44'h51422363964;
assign testcases[665] = 44'h63202142854;
assign testcases[666] = 44'h5240127199c;
assign testcases[667] = 44'h51422363964;
assign testcases[668] = 44'h41202262945;
assign testcases[669] = 44'h43532373773;
assign testcases[670] = 44'h65322273663;
assign testcases[671] = 44'h43301131879;
assign testcases[672] = 44'h54331252a5c;
assign testcases[673] = 44'h44301142987;
assign testcases[674] = 44'h44522373574;
assign testcases[675] = 44'h43222273733;
assign testcases[676] = 44'h33232383743;
assign testcases[677] = 44'h34411131a4a;
assign testcases[678] = 44'h34411131a4a;
assign testcases[679] = 44'h34411131a4a;
assign testcases[680] = 44'h43102362735;
assign testcases[681] = 44'h54702162554;
assign testcases[682] = 44'h33232263844;
assign testcases[683] = 44'h4331b362654;
assign testcases[684] = 44'h76302362548;
assign testcases[685] = 44'h44332373843;
assign testcases[686] = 44'h52312142867;
assign testcases[687] = 44'h5933d173583;
assign testcases[688] = 44'h53322383653;
assign testcases[689] = 44'h41401242877;
assign testcases[690] = 44'h52302152975;
assign testcases[691] = 44'h44211272775;
assign testcases[692] = 44'h34211272775;
assign testcases[693] = 44'h35111272785;
assign testcases[694] = 44'h63642384684;
assign testcases[695] = 44'h44332373744;
assign testcases[696] = 44'h42301131778;
assign testcases[697] = 44'h64531373574;
assign testcases[698] = 44'h64531373574;
assign testcases[699] = 44'h64532373574;
assign testcases[700] = 44'h75732273584;
assign testcases[701] = 44'h34201151aaf;
assign testcases[702] = 44'h45202132745;
assign testcases[703] = 44'h44301241646;
assign testcases[704] = 44'h33311141a5c;
assign testcases[705] = 44'h73411112227;
assign testcases[706] = 44'h44212382675;
assign testcases[707] = 44'h52412362678;
assign testcases[708] = 44'h62432244655;
assign testcases[709] = 44'h46202132643;
assign testcases[710] = 44'h43232363944;
assign testcases[711] = 44'h7340124165b;
assign testcases[712] = 44'h7340124165b;
assign testcases[713] = 44'h44421382945;
assign testcases[714] = 44'h35311272a57;
assign testcases[715] = 44'h42301252b96;
assign testcases[716] = 44'h65322183573;
assign testcases[717] = 44'h53442254353;
assign testcases[718] = 44'h42301252b96;
assign testcases[719] = 44'h63502242b56;
assign testcases[720] = 44'h43422363442;
assign testcases[721] = 44'h33402162b66;
assign testcases[722] = 44'h5430114195a;
assign testcases[723] = 44'h4430123184b;
assign testcases[724] = 44'h63401141637;
assign testcases[725] = 44'h45202252646;
assign testcases[726] = 44'h4331124198a;
assign testcases[727] = 44'h52322133474;
assign testcases[728] = 44'h41312252956;
assign testcases[729] = 44'h34308172674;
assign testcases[730] = 44'h42332153966;
assign testcases[731] = 44'h43522493854;
assign testcases[732] = 44'h83411112428;
assign testcases[733] = 44'h43332263453;
assign testcases[734] = 44'h55221173873;
assign testcases[735] = 44'h43311142654;
assign testcases[736] = 44'h43332263453;
assign testcases[737] = 44'h55221173873;
assign testcases[738] = 44'h52311252737;
assign testcases[739] = 44'h43311142654;
assign testcases[740] = 44'h5541100193c;
assign testcases[741] = 44'h32301121a68;
assign testcases[742] = 44'h52401152876;
assign testcases[743] = 44'h33231253944;
assign testcases[744] = 44'h65322163745;
assign testcases[745] = 44'h62f0124186b;
assign testcases[746] = 44'h52321293766;
assign testcases[747] = 44'h53421362529;
assign testcases[748] = 44'h52422263865;
assign testcases[749] = 44'h53421362529;
assign testcases[750] = 44'h53421362529;
assign testcases[751] = 44'h52521463666;
assign testcases[752] = 44'h42431564654;
assign testcases[753] = 44'h52321293766;
assign testcases[754] = 44'h34505152553;
assign testcases[755] = 44'h5340124185b;
assign testcases[756] = 44'h33332263a44;
assign testcases[757] = 44'h52442464ac3;
assign testcases[758] = 44'h514023528e5;
assign testcases[759] = 44'h514023528e5;
assign testcases[760] = 44'h52422263865;
assign testcases[761] = 44'h52422263865;
assign testcases[762] = 44'h53552394462;
assign testcases[763] = 44'h26041244976;
assign testcases[764] = 44'h43312262794;
assign testcases[765] = 44'h53402252348;
assign testcases[766] = 44'h47633494543;
assign testcases[767] = 44'h52301011777;
assign testcases[768] = 44'h40322243a33;
assign testcases[769] = 44'h40322243a33;
assign testcases[770] = 44'h51312242a45;
assign testcases[771] = 44'h41506352633;
assign testcases[772] = 44'h42606352633;
assign testcases[773] = 44'h43341364a44;
assign testcases[774] = 44'h83421143746;
assign testcases[775] = 44'h4250524187b;
assign testcases[776] = 44'h71401132468;
assign testcases[777] = 44'h52232374663;
assign testcases[778] = 44'h524423649b4;
assign testcases[779] = 44'h714322548a2;
assign testcases[780] = 44'h35002021938;
assign testcases[781] = 44'h63222283573;
assign testcases[782] = 44'h524423649b4;
assign testcases[783] = 44'h714322548a2;
assign testcases[784] = 44'h52232374663;
assign testcases[785] = 44'h63321243813;
assign testcases[786] = 44'h64331243813;
assign testcases[787] = 44'h64331243813;
assign testcases[788] = 44'h34221142b45;
assign testcases[789] = 44'h63321243813;
assign testcases[790] = 44'h64331243813;
assign testcases[791] = 44'h33301132a97;
assign testcases[792] = 44'h46112252665;
assign testcases[793] = 44'h33301132a97;
assign testcases[794] = 44'h64302262563;
assign testcases[795] = 44'h54322253543;
assign testcases[796] = 44'h65222283473;
assign testcases[797] = 44'h533323538a4;
assign testcases[798] = 44'h22212242a34;
assign testcases[799] = 44'h32301121978;
assign testcases[800] = 44'h63631263542;
assign testcases[801] = 44'h33522383753;
assign testcases[802] = 44'h55332383563;
assign testcases[803] = 44'h42331263a45;
assign testcases[804] = 44'h54311142745;
assign testcases[805] = 44'h63631263542;
assign testcases[806] = 44'h44332373744;
assign testcases[807] = 44'h43332373644;
assign testcases[808] = 44'h35232493633;
assign testcases[809] = 44'h43332373744;
assign testcases[810] = 44'h33522383753;
assign testcases[811] = 44'h35003142763;
assign testcases[812] = 44'h44302062a53;
assign testcases[813] = 44'h43342264a44;
assign testcases[814] = 44'h64243283576;
assign testcases[815] = 44'h43211142443;
assign testcases[816] = 44'h7241103266a;
assign testcases[817] = 44'h48221153753;
assign testcases[818] = 44'h43211142443;
assign testcases[819] = 44'h48221153753;
assign testcases[820] = 44'h44301131a7b;
assign testcases[821] = 44'h59223183373;
assign testcases[822] = 44'h52212242844;
assign testcases[823] = 44'h42212242944;
assign testcases[824] = 44'h7241103266a;
assign testcases[825] = 44'h52422263865;
assign testcases[826] = 44'h53422153976;
assign testcases[827] = 44'h6330115185c;
assign testcases[828] = 44'h51322133647;
assign testcases[829] = 44'h51302132648;
assign testcases[830] = 44'h52302243f96;
assign testcases[831] = 44'h61411262579;
assign testcases[832] = 44'h5331224196c;
assign testcases[833] = 44'h5330113174b;
assign testcases[834] = 44'h52302243f96;
assign testcases[835] = 44'h6531124164c;
assign testcases[836] = 44'h5330126183a;
assign testcases[837] = 44'h5330126183a;
assign testcases[838] = 44'h5330126183a;
assign testcases[839] = 44'h6431114263a;
assign testcases[840] = 44'h6431114263a;
assign testcases[841] = 44'h82332264652;
assign testcases[842] = 44'h82332264652;
assign testcases[843] = 44'h52301232767;
assign testcases[844] = 44'h52301241858;
assign testcases[845] = 44'h52301241858;
assign testcases[846] = 44'h42441353433;
assign testcases[847] = 44'h84301122537;
assign testcases[848] = 44'h82332264652;
assign testcases[849] = 44'h32201241959;
assign testcases[850] = 44'h52301232767;
assign testcases[851] = 44'h75532364664;
assign testcases[852] = 44'h523012428e4;
assign testcases[853] = 44'h64631253552;
assign testcases[854] = 44'h523012428e4;
assign testcases[855] = 44'h62301242ba6;
assign testcases[856] = 44'h75532364664;
assign testcases[857] = 44'h75532364664;
assign testcases[858] = 44'h42421353765;
assign testcases[859] = 44'h43318362754;
assign testcases[860] = 44'h73301232786;
assign testcases[861] = 44'h534323648a3;
assign testcases[862] = 44'h24011262975;
assign testcases[863] = 44'h4330114185b;
assign testcases[864] = 44'h24011262975;
assign testcases[865] = 44'h4330114061c;
assign testcases[866] = 44'h523012428e4;
assign testcases[867] = 44'h624322548a1;
assign testcases[868] = 44'h534313648b3;
assign testcases[869] = 44'h53301232795;
assign testcases[870] = 44'h36623163554;
assign testcases[871] = 44'h64631253552;
assign testcases[872] = 44'h43211141527;
assign testcases[873] = 44'ha1501012214;
assign testcases[874] = 44'h61301022935;
assign testcases[875] = 44'h52301152775;
assign testcases[876] = 44'h5431034183c;
assign testcases[877] = 44'h33305242736;
assign testcases[878] = 44'h41506242732;
assign testcases[879] = 44'h51301141aba;
assign testcases[880] = 44'h52301152775;
assign testcases[881] = 44'h84401043755;
assign testcases[882] = 44'h63411142669;
assign testcases[883] = 44'h63411142669;
assign testcases[884] = 44'h52331283965;
assign testcases[885] = 44'h44301141a8b;
assign testcases[886] = 44'h53301261759;
assign testcases[887] = 44'h43302231998;
assign testcases[888] = 44'h53301261759;
assign testcases[889] = 44'h43302231998;
assign testcases[890] = 44'h24012262885;
assign testcases[891] = 44'h33201241a38;
assign testcases[892] = 44'h33301242d54;
assign testcases[893] = 44'h5430124163b;
assign testcases[894] = 44'h33201241a38;
assign testcases[895] = 44'h32402121766;
assign testcases[896] = 44'h52322392766;
assign testcases[897] = 44'h53302132546;
assign testcases[898] = 44'h43301121557;
assign testcases[899] = 44'h52322392766;
assign testcases[900] = 44'h42422252968;
assign testcases[901] = 44'h63332143834;
assign testcases[902] = 44'h43332383532;
assign testcases[903] = 44'h34322372734;
assign testcases[904] = 44'h52302362452;
assign testcases[905] = 44'h72402032588;
assign testcases[906] = 44'h73402022576;
assign testcases[907] = 44'h5340124184b;
assign testcases[908] = 44'h62422163955;
assign testcases[909] = 44'h63332284562;
assign testcases[910] = 44'h44211152685;
assign testcases[911] = 44'h44212152685;
assign testcases[912] = 44'h44212152685;
assign testcases[913] = 44'h33001112923;
assign testcases[914] = 44'h64302132834;
assign testcases[915] = 44'h33001112923;
assign testcases[916] = 44'h61412252966;
assign testcases[917] = 44'h63301141328;
assign testcases[918] = 44'h5330114153a;
assign testcases[919] = 44'h72401142326;
assign testcases[920] = 44'h50312353c44;
assign testcases[921] = 44'h64621353642;
assign testcases[922] = 44'h64621353642;
assign testcases[923] = 44'h43332483745;
assign testcases[924] = 44'h63402352b57;
assign testcases[925] = 44'h43212132845;
assign testcases[926] = 44'h28112132933;
assign testcases[927] = 44'h43312362454;
assign testcases[928] = 44'h43332363d55;
assign testcases[929] = 44'h44642243653;
assign testcases[930] = 44'h6151013263a;
assign testcases[931] = 44'h43431383532;
assign testcases[932] = 44'h43332483745;
assign testcases[933] = 44'h33321372844;
assign testcases[934] = 44'h43431383532;
assign testcases[935] = 44'h43412382632;
assign testcases[936] = 44'h45302022549;
assign testcases[937] = 44'h44642243653;
assign testcases[938] = 44'h44322393965;
assign testcases[939] = 44'h63342273554;
assign testcases[940] = 44'h44321272674;
assign testcases[941] = 44'h43431383864;
assign testcases[942] = 44'h25201132c45;
assign testcases[943] = 44'h5631125163b;
assign testcases[944] = 44'h42322153842;
assign testcases[945] = 44'h41312142c46;
assign testcases[946] = 44'h74a42374344;
assign testcases[947] = 44'h71301152335;
assign testcases[948] = 44'h5a212023964;
assign testcases[949] = 44'h53411032749;
assign testcases[950] = 44'h64302152534;
assign testcases[951] = 44'h62321153555;
assign testcases[952] = 44'h41301132765;
assign testcases[953] = 44'h72402242435;
assign testcases[954] = 44'h62321153555;
assign testcases[955] = 44'h64302152534;
assign testcases[956] = 44'h64302152534;
assign testcases[957] = 44'h42302132a66;
assign testcases[958] = 44'h42301132a66;
assign testcases[959] = 44'h53342263543;
assign testcases[960] = 44'h53342263543;
assign testcases[961] = 44'h6531123267b;
assign testcases[962] = 44'h53342263543;
assign testcases[963] = 44'h42211142959;
assign testcases[964] = 44'h33231253844;
assign testcases[965] = 44'h72411132639;
assign testcases[966] = 44'h44302272634;
assign testcases[967] = 44'h52341254843;
assign testcases[968] = 44'h4030113199a;
assign testcases[969] = 44'h35100121959;
assign testcases[970] = 44'h25000131a3b;
assign testcases[971] = 44'h3320114195c;
assign testcases[972] = 44'h52341254843;
assign testcases[973] = 44'h4030113199a;
assign testcases[974] = 44'h514021429da;
assign testcases[975] = 44'h63212143653;
assign testcases[976] = 44'h41312352b46;
assign testcases[977] = 44'h41322373852;
assign testcases[978] = 44'h63311252a77;
assign testcases[979] = 44'h32707022655;
assign testcases[980] = 44'h32707022645;
assign testcases[981] = 44'h63311252a77;
assign testcases[982] = 44'h25201121b4c;
assign testcases[983] = 44'h34311131a4a;
assign testcases[984] = 44'h52302352a67;
assign testcases[985] = 44'h35202242a66;
assign testcases[986] = 44'h63312262656;
assign testcases[987] = 44'h63312262646;
assign testcases[988] = 44'h52302352a67;
assign testcases[989] = 44'h6342104253a;
assign testcases[990] = 44'h71411252336;
assign testcases[991] = 44'h73402022676;
assign testcases[992] = 44'h43342483735;
assign testcases[993] = 44'h53202022a55;
assign testcases[994] = 44'h72301173864;
assign testcases[995] = 44'h63302152546;
assign testcases[996] = 44'h33302012886;
assign testcases[997] = 44'h43323253954;
assign testcases[998] = 44'h63342264553;
assign testcases[999] = 44'h62602362565;


  
  localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
  wire [$clog2(CLASS_CNT)-1:0] prediction;

  // Instantiate module under test
 winequality_white_bs #() dut (
    .features(sample),
    .clk(clk),
    .rst(rst),
    .prediction(prediction)
  );
  
  always #halfPeriod clk <= ~clk;

  integer i;
  initial begin
    $write("["); //"
    for(i=0;i<TEST_CNT;i=i+1)
        runtestcase(i);
    $display("]");
    $finish;
  end

  localparam [$clog2(CLASS_CNT)-1:0] maxclass = CLASS_CNT-1;

  task runtestcase(input integer i); begin
    sample <= testcases[i];
    rst <= 1;
    clk <= 0;
    #period
    rst <= 0;
    #period
    #((FEAT_CNT+HIDDEN_CNT-1)*period)
    $write("%d, ",(maxclass-prediction));
  end
  endtask

endmodule
