
















module cardio_bnn1_bnnpaarter #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 8880'h001500aa0001001400a90001001500a70001005400a50001001e00a40001001400a10001002e009f00010042009e0001002a009d00010090009c0001002f009b00010052009a0001003f00990001003b00970001005c00950001004800940001002100920001001e008f0001005b008e00010058008d00010026008c0001002e008b0001002600870001004000860001007600850001003a00840001005a00830001006e00820001006f008100010079008000010037007f00010046006d0001005800590001003e00960000006700930000006b00910000007b008a00000060008900000049007e00000048007d0000006a007c0000006c007a0000004700780000006500770000005d00750000004c00740000006300730000005500720000003e00710000003400700000005e00690000005600680000005900660000002f00640000003d006200000046006100000031005f00000051005b00000041005a0000002b00570000003a00560000002d00550000004000540000005100530000004300530000004b00500000003700500000004d004f00000045004f0000004c004e0000003d004e00000034004d00000040004b0000004400490000003500470000004100450000002f00440000002200430000003900420000003100420000002800410000003d003f0000002e003f00000033003e0000002c003c0000001500390000003500380000001a00380000003400360000001400360000001e00350000002c00330000002700300000001800300000002e002f0000002c002d00000025002c00000029002b00000026002b0000001e002a0000001b002a0000002700290000001e00290000001800290000001a00270000002500260000001400260000001b00310001001800300001001a00270001001400570000003300520000001b003700000024004a00010036003800010021003500010008003200010026002f00010015002a0001001c002300010022003c00000014003b00000025003a0000002700390000002900340000002d003000000021002e0000001900240000001d00230000002000210000001f00210000001a001f0000002b00310001001e002900010027002800010025003300000015002900000027002c0001001b002200010025002b00000025002a00000016001c00000018001f0000001f002d0001000800320000001700200001002000240000001b001e0000001800260001001d00230001001700200000001b001e00010019002400010001000300010015001a0000001c00230000001f002100010016001d00010014002800000016001d0000001b002200000017001900000017001900010008001300010009001000000016001c00010005000a00010000000c00010004000f00000002001100000014001a00000006000d0000000e001200000015001800000007000b00000007000b0001000e001200010008001300000006000d00010002001100010000000c00000004000f00010005000a0000000900100001000100030000 ;
localparam YMAP = 1280'h000000b3000100cb000000c2000000a8000100c5000000c4000100bc000100b2000100b0000000ca000000b1000100b8000100af000000b9000000c8000100be000000c7000000ac000100ad000000a6000000c3000100b4000100ab000100b6000000c6000000bf000000a2000000c1000000ae000000c9000000a000010098000000bd000000b7000000c000010088000000ba000000a3000100b5000000bb;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 120'b101010000001111100000011001000100011100111001011000110110011011101101001101001110100101100111001001101110110000110110011 ;
localparam WIDTH = 320'h08070708080808080708070707080707060807080707070707070808080807080707070707070708;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;
generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam subad = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(subad)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] < 0;
    initial begin
        #20
        $display("%b, %d | %d", signy, ymap, node[ymap]);
    end
end
endgenerate

initial begin
    #10
    for(j=0;j<FULLCNT;j=j+1) begin
        $display("%d | %d | %b, %d, %d", j, node[j], PAAR0[(j- FEAT_CNT )*48],  PAAR0[(j-FEAT_CNT)*48+16+:16], PAAR0[(j-FEAT_CNT)*48+32+:16]);
    end
end

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wneur[j])
            tmpscore = tmpscore + hidden[j];
        else 
            tmpscore = tmpscore + hidden_n[j];
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = tmpscore;
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
