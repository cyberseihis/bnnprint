module tst ();

wire out1;
wire out2;

compare1side c1 (
31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd73741824, 31'd73741824, 31'd73741824, 31'd73741824, 31'd73741824,
out1);

compare2side c2 (
31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd12, 31'd73741824, 31'd73741824, 31'd73741824, 31'd73741824, 31'd73741824,
out2);

initial begin
    #1
    $display("c1 %b",out1);
    $display("c2 %b",out2);
end

endmodule
