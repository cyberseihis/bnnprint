`timescale 1us/1ns









module tbgasId_tnn1_tnnpar #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)();
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
reg clk;
reg [FEAT_CNT*FEAT_BITS-1:0] features;
wire [$clog2(CLASS_CNT)-1:0] prediction;
wire [FEAT_CNT*FEAT_BITS-1:0] testcases [TEST_CNT-1:0];
parameter Nsperiod=5000;
localparam period=Nsperiod/500;


assign testcases[0] = 512'hfef00012fef00012fff00112fff00012fff00012fff00012fff00001fff00001fef00003fef00003fff00003fff00002fff00005fff00014fff00001fef00001;
assign testcases[1] = 512'hfef00012fef00012fff00122fff00122fef00012fef00112fff01101fff00101fef00004fef00003fff00003fff00002fff00005fff00014fff00101fef00101;
assign testcases[2] = 512'hfef00122fef00122ffe00123ffe00123fef00123fef01113fef11101fff01101fef00104fef00104ffe00004fff00003fff00005fff00015fff00102fef01101;
assign testcases[3] = 512'hfef00122fef01122ffe00223ffe00223fef01123fef01113fef11101fff11101fef00104fef00104ffe00004fff00003fff00005fff00115fff01102fef11101;
assign testcases[4] = 512'hfef00123fef01122ffd00234ffe00233fef01123fef01123fee11102fee11102fef00104fef00104ffe00004fff00003fff00015fff00125ffe01102fef01102;
assign testcases[5] = 512'hfdf10133fdf01133ffc01344ffd01244fee01133fee01223fde12212fee12212fde00105fde00105ffd00105fff00104fff00016ffe00125fee01203fde02202;
assign testcases[6] = 512'hfde10233fde01233ffb01345ffc01345fee01234fee11224fdd23213fed12213fde01105fde01205ffc00106fff00105fff00016ffe00136fed01203fde12203;
assign testcases[7] = 512'hfde10244fde01244feb01455ffc01355fde01244fde11234fdd23313fdd13313fde01205fde01205ffb00106fff00105fff00016fed00136fed02303fdd13203;
assign testcases[8] = 512'hfcd10254fde12254fea01466feb01366fdd02244fdd12234edc23313fdd23313fdd01206fdd01206ffb00107fff00106fff00017fed00146fed02304fdd13303;
assign testcases[9] = 512'hfcd10354fcd12254fe901467fea01366fdd02255fdd12335ecc24314fdc23314fcd11206fcd01206fea00107ffe00106fff00017fec00147fec02304fdd13303;
assign testcases[10] = 512'hfcd11365fcd12365fe801477fe901477fcc12355fcc12345ecc24414fdc24314fcc11206fcc01206fe900108ffe00107ffe00017fec00147fec02404ecd14304;
assign testcases[11] = 512'hfbc11365fcc12365fe701578fe901477fcc12355fcc12346ecc34414fdc24414fcc11207fcc11207fe800108ffe00107ffe00018feb00157fec03405fcc14304;
assign testcases[12] = 512'hfbc11365fbc12365fe601588fe801488fcb12366fcb12346ecb35415edb24414fcb11207fbb11307fe800109ffe00107ffe00018feb00258fec03405ecc15404;
assign testcases[13] = 512'hfbb11375fbb12376fe601588fe701488fcb12366fbb12356ecb35415fdb25415fbb11307fbb11307fe700109ffe00108ffe00018fda00258fdb03405ecc15404;
assign testcases[14] = 512'hfef00012fef00012fff00112fff00112fff00012fff00012fff00001fff00001fef00003fef00003fff00003fff00002fff00005fff00014fff00001fef00001;
assign testcases[15] = 512'hfef00112fef00112ffe00123fff00123fef00113fef00113fef01101fff01101fef00004fef00104fff00003fff00003fff00005fff00015fff00101fef01101;
assign testcases[16] = 512'hfef00122fef01122ffe00223ffe00123fef01123fef01113fef11101fff01101fef00104fef00104ffe00004fff00003fff00005fff00015fff01102fef01101;
assign testcases[17] = 512'hfef00123fef01123ffd01234ffe00233fef01123fef01113fee11102fff11102fef00104fef00104ffe00004fff00004fff00005fff00125ffe01102fef01102;
assign testcases[18] = 512'hfdf00123fef01123ffd01334ffd01234fef01123fef01213fee12212fee12202fef00104fef00104ffd00105fff00104fff00006ffe00125ffe01202fef01102;
assign testcases[19] = 512'hfde10233fde01233ffc01345ffc01344fee01234fee11224fde12212fee12212fde01105fde01205ffc00105fff00105fff00016ffe00126fee01203fde02202;
assign testcases[20] = 512'hfde10234fde02234feb01446ffc01345fde01234fde12224edd23313fed13213fde01205fdd01205ffb00106fff00105fff00016fed00136fed02303fde12203;
assign testcases[21] = 512'hfcd11344fdd12244fea01456feb01456fdd02234fdd12335fdd23313fed13313fdd11206fcd01206ffb00107fff00106fff00017fed00137fed02303fdd13303;
assign testcases[22] = 512'hfcd11344fcd12344fe901467fea01466fdd12345fdd12335edc23313fdd13313fcd11206fcd01206fea00107ffe00106ffe00017fec00137fed02304fdd13303;
assign testcases[23] = 512'hfcd11355fcd12355fe801567fea01467fcc12345fcc12335ecc24314fdc24314fcc11207fcc11306fe900108ffe00107ffe00017fec00147fec02304fdd13303;
assign testcases[24] = 512'hfbc11355fcc12355fe701568fe901477fcc12355fcc12446ecc24414fdc24414fcc11307fbc11307fe900108ffe00107ffe00018feb00248fec02404fcd14304;
assign testcases[25] = 512'hfbc11465fbc12365fe602578fe801578fcb12356fcb12446ecc34414fdc24414fbb11307fbb11307fe701109ffe00108ffe00018fea00258fec02404fcd14304;
assign testcases[26] = 512'hfbb11466fbb12466fe602679fe701578fbb13466fbb13446ecb35415fdc24414fbb11307fbb11307fe701109ffd01108ffe00118fda00258fec03405fcc14404;
assign testcases[27] = 512'hfab11476fab12476fd502689fe701588fba13466fba13457ecb35415fdb24415fba11308faa11308fe60110affd01108ffd00119fda00259fdb03405ecc15404;
assign testcases[28] = 512'hfef00012fef00012fff00112fff00012fff00012fff00012fff00001fff00001fef00003fef00003fff00003fff00002fff00005fff00014fff00001fef00001;
assign testcases[29] = 512'hfef00112fef00012ffe00123fff00122fef00112fef00112fef01101fff01101fef00004fef00004fff00003fff00003fff00005fff00015fff00101fef01101;
assign testcases[30] = 512'hfef00122fef01122ffe00223ffe00123fef01113fef01113fef11101fff01101fef00104fef00104ffe00004fff00003fff00005fff00015fff01102fef01101;
assign testcases[31] = 512'hfef00122fef01122ffd00234ffe00233fef01123fef01113fee11102fff11102fef00104fef00104ffe00004fff00003fff00005fff00125ffe01102fef01102;
assign testcases[32] = 512'hfdf00123fef01123ffd01334ffd01234fef01123fef01123fee12202fee12202fef00104fef00104ffd00104fff00104fff00016fff00125ffe01202fef01102;
assign testcases[33] = 512'hfde10233fde01233ffc01345ffd01344fee01234fee01224fde12212fee12212fde00105fde00105ffc00105fff00104fff00016ffe00136fee01203fde02202;
assign testcases[34] = 512'hfde10243fde01243ffb01455ffc01355fde01234fde11224fdd23313fed13213fde01205fde01205ffc00106fff00105fff00016ffe00136fed02303fde12203;
assign testcases[35] = 512'hfde10254fde01254fea01456ffb01355fdd01244fdd12234fdd23313fed13313fdd01206fdd01206ffb00106fff00105fff00017fed00146fed02303fdd13203;
assign testcases[36] = 512'hfcd11354fcd12354fea01566feb01466fdd12345fdd22335edc24313fdd24313fcd11206fcd01206ffa00107ffe00106fff00017fed00147fed02304fdd14303;
assign testcases[37] = 512'hfcd11355fcd12355fe901467fea01466fdc12355fcc12335ecc24314fdc24314fcc11206fcc01206fe900108ffe00106ffe00017fec00147fec02304fdd13303;
assign testcases[38] = 512'hfbc11365fcc12365fe801577fe901477fcc12355fcc12346ecc24414fdc24414fcc11207fcc11307fe900108ffe00107ffe00018feb00247fec02404fcd14304;
assign testcases[39] = 512'hfbc11365fbc12365fe701578fe901477fcc12366fcc12346ebb34414edc24414fcc11207fbb11307fe800108ffe00107ffe00018feb00258fdc03405ecc14304;
assign testcases[40] = 512'hfbc11475fbb12375fe601588fe801488fcb12366fcb12456ecb35415fdc24414fbb11307fbb11307fe700109ffe00108ffe00018fda00258fec03405ecc14404;
assign testcases[41] = 512'hfab11476fab12476fe602689fe701588fcb12466fbb13456ecb35415fdb25415fbb11307fbb11308fe701109ffe00108ffe00118fda00258fdb03405ecc15404;
assign testcases[42] = 512'hfef00012fef00012fff00112fff00012fff00012fff00012fff00001fff00001fef00003fef00003fff00003fff00002fff00005fff00014fff00001fef00001;
assign testcases[43] = 512'hfef00112fef00012fff00123fff00122fef00012fef00112fef01101fff01101fef00004fef00004fff00003fff00003fff00005fff00015fff00101fef01101;
assign testcases[44] = 512'hfef00122fef01122ffe00223ffe00123fef01123fef01113fef11101fff01101fef00104fef00104ffe00004fff00003fff00005fff00015fff01102fef01101;
assign testcases[45] = 512'hfef00122fef01122ffe00233ffe00233fef01123fef01113fef11101fff11101fef00104fef00104ffe00004fff00003fff00005fff00115fff01102fef01101;
assign testcases[46] = 512'hfef00123fef01122ffd01234ffe00233fef01123fef01113fee12212fee11102fef00104fef00104ffd00105fff00004fff00005fff00125ffe01102fef01102;
assign testcases[47] = 512'hfdf10233fdf01133ffc01344ffd01344fee01233fee11223fdd12212fee12212fde01105fde01205ffd00105fff00104fff00016ffe00126fee01203fde02202;
assign testcases[48] = 512'hfde10233fde01233ffb01455ffc01355fee01234fee11224fdd23313fed13313fde01205fde01205ffc00106fff00105fff00016ffe00136fed02303fde13203;
assign testcases[49] = 512'hfde10244fde12244feb01456ffc01355fde01234fde12234fdd23313fed13313fdd01206fdd01206ffb00106fff00105fff00017fed00136fed02303fde13303;
assign testcases[50] = 512'hfcd11244fce12244fea01466feb01366fdd02244fdd12234ecc24414fdc24314fcd11206fcd01206ffa00107ffe00106fff00017fed00137fed02304fdd13303;
assign testcases[51] = 512'hfcd11354fcd12254fe901467fea01466fdd12245fdd12335ecc24414fdc24414fcc11206fcc01206fea00107ffe00106ffe00017fec00147fec02304fdd13303;
assign testcases[52] = 512'hfcd11355fcd12355fe801567fe901477fcc12355fcc12345ecc24414fdc24414fcc11207fcc11307fe900108ffe00107ffe00018feb00247fec02404fdd13304;
assign testcases[53] = 512'hfbc11365fcc12365fe801578fe901477fcc12355fcc12345ecb34415fdc24414fbb11307fbb11307fe800109ffe00107ffe00018feb00258fec02404fcd14304;
assign testcases[54] = 512'hfbc11365fbc12365fe701578fe801487fcc12365fcc12346ecb35415fdb25415fbb11307fbb11307fe700109ffe00108ffe00018fea00258fec03405ecc14404;
assign testcases[55] = 512'hfbb11365fbb12375fe601588fe701488fcb12366fbb12346ecb35515fdb25415fba11308fba11308fe70110affd00108ffd00019fda00259fec03405ecc14404;
assign testcases[56] = 512'hfef00012fef00012fff00022fff00012fff00012fff00012fff00001fff00001fef00003fef00003fff00003fff00002fff00005fff00014fff00001fef00001;
assign testcases[57] = 512'hfef00122fef00112ffe00123fff00122fef00112fef00112fef01101fff01101fef00004fef00104fff00003fff00003fff00005fff00015fff00101fef01101;
assign testcases[58] = 512'hfef00122fef01122ffe00233ffe00133fef01123fef01113fef11101fff01101fef00104fef00104ffe00004fff00003fff00005fff00025fff01102fef01101;
assign testcases[59] = 512'hfef00123fef01123ffd00234ffe00233fef01123fef01123fee11112fee11102fef00104fef00104ffe00004fff00004fff00016fff00125ffe01102fef01102;
assign testcases[60] = 512'hfdf10123fdf01123ffd01334ffd01234fef01123fef01123fee12212fee12212fef00105fde00105ffd00105fff00104fff00016ffe00125ffe01202fef01102;
assign testcases[61] = 512'hfde10233fde01233ffc01345ffd01344fee01234fee11224fdd12213fee12212fde01105fde01205ffc00105fff00105fff00016ffe00136fee01203fde02202;
assign testcases[62] = 512'hfde10233fde01243ffb01455ffc01355fee01234fde12224fdd23313fed13313fde01205fde01205ffc00106fff00105fff00016fed00136fed02303fde12203;
assign testcases[63] = 512'hfde11244fde12244fea01456ffb01455fde02244fde12234fdd24313fed23313fdd11206fdd01206ffb00107fff00106fff00017fed00136fed02303fdd13303;
assign testcases[64] = 512'hfcd11354fcd12254fea01466feb01466fdd02244fdd12335ecc24414fdc24314fcd11206fcd01206ffa00107ffe00106fff00017fec00147fed02304fdd13303;
assign testcases[65] = 512'hfcd11354fcd12354fe901467fea01466fdd12355fdd12345ecc24414fdc24414fcc11206fcc01306fea00108ffe00106ffe00017fec00147fec02304fdd13304;
assign testcases[66] = 512'hfcd11355fcd12365fe801577fe901477fcc12355fcc12345ecc24414fdc24414fcc11207fcc11307fe900108ffe00107ffe00018feb00247fec02404fdd14304;
assign testcases[67] = 512'hfbc11365fcc12365fe801578fe901477fcc12355fcc12345ecb35415fdc24414fbb11307fbb11307fe800108ffe00107ffe00018feb00258fec02404fcd14304;
assign testcases[68] = 512'hfbc11365fbc12375fe701588fe801488fcc12366fcc12346ecb35415edb25415fbb11307fbb11307fe800109ffe00108ffe00018fea00258fec03405ecc14404;
assign testcases[69] = 512'hfbb11475fbb12375fe601588fe801488fcb12366fcb12356ecb35515fdb25415fba11308fba11308fe701109ffe00108ffe00019fda00258fec03405ecc14404;
assign testcases[70] = 512'hfef00012fef00012fff00112fff00012fff00012fff00012fff00001fff00001fef00003fef00003fff00003fff00002fff00005fff00014fff00001fef00001;
assign testcases[71] = 512'hfef00112fef00112ffe00123fff00123fef00112fef00112fef01101fff01101fef00004fef00104fff00003fff00003fff00005fff00015fff00101fef01101;
assign testcases[72] = 512'hfef00112fef01112ffe00223ffe00123fef01113fef01113fef11101fff01101fef00104fef00104ffe00004fff00003fff00005fff00015fff01102fef01101;
assign testcases[73] = 512'hfef00123fef01122ffd01234ffe00233fef01123fef01113fee11102fee11102fef00104fef00104ffe00104fff00004fff00005fff00125fff01102fef01102;
assign testcases[74] = 512'hfdf00223fdf11123ffd01334ffd01234fef11223fef12213fee44212fee34212fef11105fdf11205ffd00105fff00104fff00006ffe00125ffe12202fef13202;
assign testcases[75] = 512'hfde10223fde01223ffc01345ffd01344fee01224fee11224fdd12213fee12212fde01105fde01205ffc00106fff00105fff00016ffe00126fee01203fde02202;
assign testcases[76] = 512'hfde10234fde12234ffb01445ffc01345fde02234fde12224edd23313fed13313fdd01206fdd01206ffb00106fff00105fff00017fed00126fed02303fde12203;
assign testcases[77] = 512'hfce11334fde12234fea01456feb01456fdd02234fdd12324fdd23313fed13313fcd11206fcd01206ffb00107fff00106fff00017fed00137fed02303fde13303;
assign testcases[78] = 512'hfcd11344fcd12344fe901557fea01466fdd12345fdd12335ecc24414fdc23314fcc11206fcc01306fea00108ffe00106ffe00017fec00137fed02304fdd13303;
assign testcases[79] = 512'hfcd11355fcd12355fe901567fea01467fdc12345fcc12335ecc24414fdc24414fcc11307fcc11307fe900108ffe00107ffe00018feb00248fed02304fdd13303;
assign testcases[80] = 512'hfbc11355fbc12355fe801567fe901477fcc12355fcc12345ecc24414fdc24414fbb11307fbb11307fe800108ffe00107ffe00018feb00248fec02404fdd14304;
assign testcases[81] = 512'hfbc11465fbc12365fe702578fe801477fcc12355fcc12346ecb34415fdc24414fbb11307fbb11308fe801109ffe00108ffe00018fea00258fec02404fdd14304;
assign testcases[82] = 512'hfbc11465fbb12465fe602578fe801588fcb12366fcb12446ecb35415fdb24415fba11308fba11308fe701109ffe00108ffd00119fda00259fec03405fcd14404;
assign testcases[83] = 512'hfbb11476fbb12476fe602689fe801588fcb12366fbb12456ecb35515fdb25415fba11308fba11408fe70110affe00108ffd00129fda00269fec03405fcc14404;
assign testcases[84] = 512'hfef00012fef00012fff00012fff00012fff00012fef00012fff00000fff00000fef00004fef00003fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[85] = 512'hfde00233fde01233ffd00233ffe00233fee01233fde01224fff00000fff00000fde00105fde00105ffd00004fff00003fff00016fee00136fff00001fef00001;
assign testcases[86] = 512'hfef11301fef12301fff01401fff01301fff12302fff13402fff00000fff00000fef11303fef01303fff00102fff00101fff00104fff00204fff00000fff00000;
assign testcases[87] = 512'hfde11344fcd12344ffc01344ffd01344fdd12344fdd12335fff00000fff00001fdd11206fdd01306ffc00105fff00104ffe00017fec00247fff00001fef00001;
assign testcases[88] = 512'hfbc11475fbc13475fe901466fea01365fcb13476fba14567fff00000fff00101fbb11307fbb12407fea00107ffe00106ffd00129fd901369fff00001fef00001;
assign testcases[89] = 512'hfbb21586fab14596fe801577fea01466fba13587fa924678fff00001fff01101fba12408fba12408fe901108ffe00106ffc0012afd70137afff00001fef01001;
assign testcases[90] = 512'hfef00012fef00012fff00012fff00012fff00012fef00012fff00000fff00000fef00003fef00003fff00003fff00002fff00005fff00014fff00001fff00000;
assign testcases[91] = 512'hfdf10233fde01233ffd00233ffe00233fee01233fee11234fff00000fff00000fde00105fde01205ffe00004fff00003fff00016ffe00136fff00001fef00001;
assign testcases[92] = 512'hfde11354fdd12354ffc01344ffd01244fdd12344fdd12345fff00000fff00001fdd11206fdd01206ffc00105fff00104ffe00017fec00247fff00001fef00001;
assign testcases[93] = 512'hfcd11465fcd13465fea01455ffc01355fcc13465fcb13456fff00000fff00001fcc11307fcc11307ffb00106fff00105ffe00119fda01268fff00001fef00001;
assign testcases[94] = 512'hfbc21475fbc13486fe901466feb01366fbb13476fba14567fff00000fff00001fbb11307fbb12407fea00107ffe00106ffd00129fd901379fff00001fef00001;
assign testcases[95] = 512'hfab21586fbb14596fe801577fea01476fba14587fa924678fff00001fff01101fba12408fba12408fe901108ffe00107ffc0012afc70138afff00001fef01001;
assign testcases[96] = 512'hfef00022fef00022fff00012fff00012fff00012fef00012fff00000fff00000fef00004fef00003fff00003fff00002fff00005fff00025fff00001fff00000;
assign testcases[97] = 512'hfde00233fde01233ffd00233ffe00233fee01234fee11234fff00000fff00000fde00105fde01205ffe00104fff00003fff00016ffe00136fff00001fef00001;
assign testcases[98] = 512'hfcd11354fcd12354ffc01344ffd01344fdd12355fdc13445fff00000fff00001fdd11206fcd01306ffc00105fff00104ffe00017fec00247fff00001fef00001;
assign testcases[99] = 512'hfcd11465fcd13465feb01455ffc01355fcc13465fcb13456fff00000fff00001fcc11307fcc11307ffb00106fff00105ffe00128fda01268fff00001fef00001;
assign testcases[100] = 512'hfbc21475fbc13486fe901466ffb01366fcb13476fba24568fff00001fff01101fcb11308fbb12407ffa00107ffe00106ffd0012afd901379fff00001fef00001;
assign testcases[101] = 512'hfab21596fbb14596fe801577fea01476fba14597fa824679fff00001fff01101fba12408fba12408fe901108ffe01107ffc0012afc70138afff00101fef01001;
assign testcases[102] = 512'hfef00012fef00012fff00012fff00012fff00012fef00012fff00000fff00000fef00004fef00003fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[103] = 512'hfde00233fde01233ffd00233ffe00223fee01234fde11224fff00000fff00000fde00105fde01205ffe00104fff00003fff00016ffe00136fff00001fef00001;
assign testcases[104] = 512'hfcd11344fcd12344ffc01345ffd01344fdd12345fcc13435fff00000fff00001fcd11206fcd01306ffc00105fff00104ffe00017fec00247fff00001fef00001;
assign testcases[105] = 512'hfcd11455fcc13465fea01456ffb01355fcc13456fbb14546fff00000fff00001fcc11307fcc11307ffb00106fff00105ffe00119fda01259fff00001fef00001;
assign testcases[106] = 512'hfbc21576fbb14576fe901566fea01466fba14577fa924668fff00000fff00101fbb12408fbb12408fea00107ffe00106ffd0012afd80137afff00001fef00001;
assign testcases[107] = 512'hfab21596fab14596fe801577fe901476fb914587fa825679fff00001fff01101fba12408faa12408fe901108ffe00107ffc0012bfc70138bfff00101fef01001;
assign testcases[108] = 512'hfef00012fef00012fff00012fff00012fef00012fef00012fff00000fff00000fef00004fef00004fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[109] = 512'hfde10233fde01233ffd00233ffe00233fee01234fde12234fff00000fff00000fde01205fde01205ffe00104fff00103fff00016fee00136fff00001fef00001;
assign testcases[110] = 512'hfcd11354fcd12354ffc01345ffd01344fdd12355fcc13446fff00000fff00001fcd11306fcd11306ffc00105fff00104ffe00118fec00248fff00001fef00001;
assign testcases[111] = 512'hfcc11465fcc13465fea01456ffb01355fcc13466fbb14557fff00000fff00001fcc11307fcc11307ffb00106fff00105ffe00129fda01269fff00001fef00001;
assign testcases[112] = 512'hfbc11595fbc135a6fe901566feb01466fcb13586fba24678fff00001fff00101fbb11407fbb11407ffa00107ffe00106ffd0012afd90138afff00001fef00001;
assign testcases[113] = 512'hfab21596fab14596fe801577fe901466fba14587f9825679fff00001fff01101faa12408faa12408fe801108ffe01107ffc0012bfc70138bfff00001fef01001;
assign testcases[114] = 512'hfef00022fef00022fff00012fff00012fef00012fef00013fff00000fff00000fef00004fef00003fff00003fff00002fff00005fff00025fff00001fff00000;
assign testcases[115] = 512'hfde10233fde01243ffd00233ffe00233fee01234fde12234fff00000fff00000fde00105fde01205ffe00104fff00003fff00016ffe00136fff00001fef00001;
assign testcases[116] = 512'hfcd11354fcd12354ffc01344ffd01344fdd12355fcc13445fff00000fff00001fcd11206fcd01306ffc00105fff00104ffe00118fec00247fff00001fef00001;
assign testcases[117] = 512'hfcd11465fcc13475fea01455ffc01355fcc13466fbb14557fff00000fff00001fcc11307fcc11407ffb00106fff00105ffe00129fda01369fff00001fef00001;
assign testcases[118] = 512'hfbc21585fbb13586fe901466fea01466fbb14576fa924668fff00001fff01101fbb11307fbb12407fea00107ffe00106ffd0012afd80137afff00001fef00001;
assign testcases[119] = 512'hfab21596fab14596fe801577fea01476fba14587fa825679fff00001fff01101fba12408fba12408fe901108ffe01106ffc0012bfd70138bfff00101fef01001;
assign testcases[120] = 512'hfef00022fef00022fff00012fff00012fff00012fef00012fff00000fff00000fef00004fef00003fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[121] = 512'hfdf00233fdf01233ffe00233ffe00233fee01234fee11224fff00000fff00000fde00105fde01205ffe00004fff00003fff00016ffe00136fff00001fef00001;
assign testcases[122] = 512'hfde11344fcd12354ffc01344ffd01344fdd12345fcc13435fff00000fff00001fdd11206fdd01306ffc00105fff00104ffe00117fec00247fff00001fef00001;
assign testcases[123] = 512'hfcd11465fcc13465feb01455ffc01355fcc13455fbb14556fff00001fff00001fcc11306fcc11306ffb00106fff00105ffe00118fda01258fff00001fef00001;
assign testcases[124] = 512'hfbc11475fbc13485fea01466feb01365fcb14476fba24567fff00001fff01101fbb11307fbb12407fea00107ffe00106ffd00129fd901369fff00001fef00001;
assign testcases[125] = 512'hfbb21586fab14596fe801577fea01466fba14587fa825669fff00001fff01101fba12408fba12408fe900107ffe00106ffc0012afc70137bfff00101fef01001;
assign testcases[126] = 512'hfef00132fef01132ffe00123fff00122fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00016ffe00125fff00001fef00001;
assign testcases[127] = 512'hfde10253fde01253ffd00334ffd00233fde02244fdd12345fff00000fff00001fde01205fde01205ffd00105fff00104fff00017fed00147fff00001fef00001;
assign testcases[128] = 512'hfcd11364fcd12364ffb01445ffc01344fcc13455fcc13556fff00000fff00001fcd11306fcd11306ffc00106fff00105ffe00118feb00258fff00001fef00001;
assign testcases[129] = 512'hfcc11475fcc13475fea01456ffb01355fcb13476fba24567fff00001fff00001fcc11307fcc11307ffb00106fff00105ffd00129fd901269fff00001fef00001;
assign testcases[130] = 512'hfbb21586fbb13596fe901466fea01366fba14587fa924678fff00001fff01101fbb11308fbb12408fea00107ffe00106ffd0012afd80138afff00101fef01001;
assign testcases[131] = 512'hfef00132fef01132ffe00123fff00122fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00016ffe00125fff00001fef00001;
assign testcases[132] = 512'hfde10243fde02253ffd01334ffe00233fde02244fdd12335fff00000fff00000fde01205fde01205ffd00104fff00104fff00017fed00147fff00001fef00001;
assign testcases[133] = 512'hfcd11364fcd12364ffb01355ffc01354fdc13365fcc13456fff00000fff00001fcd11306fcd11306ffc00105fff00105ffe00118feb00258fff00001fef00001;
assign testcases[134] = 512'hfbc11475fbc13485fea01466feb01355fcb13476fba14567fff00000fff00101fbc11307fbb11307ffb00106fff00105ffd00129fd901379fff00001fef00001;
assign testcases[135] = 512'hfbb21586fbb14596fe901466fea01466fba14587fa925678fff00001fff01101fbb11408fbb12408fea00107ffe00106ffd0012afd80138afff00101fef00001;
assign testcases[136] = 512'hfef00133fef01133ffe00123fff00122fef01133fef01223fff00000fff00000fef00104fef00104ffe00003fff00003fff00016ffe00136fff00001fef00001;
assign testcases[137] = 512'hfde10244fde12244ffd01334ffd00233fdd12344fdd12335fff00000fff00001fde01205fde01205ffd00105fff00104fff00017fed00247fff00001fef00001;
assign testcases[138] = 512'hfcd11464fcd13464ffb01455ffc01344fcc13455fcb13556fff00000fff00001fcc11306fcc11306ffc00106fff00105ffe00118feb00258fff00001fef00001;
assign testcases[139] = 512'hfbc11475fbc13485fea01466ffb01355fcb13476fba24667fff00001fff00101fbb11307fbb12407ffa00107fff00106ffd00129fd901369fff00001fef00001;
assign testcases[140] = 512'hfab21586fbb14586fe801567fea01466fba14577fa825769fff00001fff01101fba12408fba12408fe901108ffe00106ffc0012afd70137afff00101fef00001;
assign testcases[141] = 512'hfaa215a7faa145b7fe701578fe901477fa915598f972578afff01101fff01101fa912409fa912409fe801109ffe01107ffc0012bfc60139bfff00101fef01001;
assign testcases[142] = 512'hfaa21597faa145a7fe702578fe901477fa915598f972578afff01001fff01101fa912409fa912509fe801108ffe01107ffc0012bfc60138bfff00101fef01001;
assign testcases[143] = 512'hfaa21596faa145a7fe701577fe901477fa915598f972578afff00001fff01101fa912409fa912509fe801108ffe01107ffc0012bfc60139bfff00101fef01001;
assign testcases[144] = 512'hfef00122fef01122ffe00223fff00122fef01123fef01223fff00000fff00000fef00104fef00104ffe00003fff00003fff00016ffe00125fff00001fef00001;
assign testcases[145] = 512'hfde10233fde02243ffd01334ffd00233fde12234fdd12335fff00000fff00001fde01205fde01205ffd00105fff00104fff00017fed00137fff00001fef00001;
assign testcases[146] = 512'hfcd11454fcd13454ffb01445ffc01344fcc13445fcb13546fff00000fff00001fcc11306fcc11306ffc00106fff00105ffe00118feb00248fff00001fef00001;
assign testcases[147] = 512'hfbc11465fbc13475fea01456feb01355fcb13466fba24557fff00001fff00101fbc11307fbb11407feb00106fff00105ffd00119fd901359fff00001fef00001;
assign testcases[148] = 512'hfbb21576fab14586fe901567fea01466fba14577fa925668fff00001fff01101fba12408fba12408fe901107ffe00106ffd0012afd80137afff00101fef00001;
assign testcases[149] = 512'hfab21597faa14597fe701578fe901477fa914588f9725779fff01001fff01101fa912408fa912409fe801108ffe01107ffc0012bfc60138bfff00101fef01001;
assign testcases[150] = 512'hfef00123fef01122ffe00223fff00122fef01123fee01223fff00000fff00000fef00104fef00104ffe00003fff00003fff00016ffe00126fff00001fef00001;
assign testcases[151] = 512'hfde11344fde12344ffc01334ffd01234fdd12344fdd13435fff00000fff00000fdd11205fdd01205ffd00105fff00104ffe00017fec00247fff00001fef00001;
assign testcases[152] = 512'hfcd11465fcd13465feb01455ffc01345fcc13455fcb14547fff00000fff00001fcc11306fcc11306ffb00106fff00105ffe00119fea01258fff00001fef00001;
assign testcases[153] = 512'hfef00012fef00022fff00012fff00012fef00012fef00013fff00000fff00000fef00004fef00004fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[154] = 512'hfde10233fde01233ffd00233ffe00233fee01234fde12334fff00000fff00000fde01105fde01205ffe00104fff00103fff00017fed00136fff00001fef00001;
assign testcases[155] = 512'hfcd11354fcd12354ffc01345ffd01344fdd13355fcc13446fff00000fff00001fcd11306fcd11306ffc00105fff00104ffe00118feb00248fff00001fef00001;
assign testcases[156] = 512'hfaa21697faa156a7fe602578fe801477f9815698f872688afff00001fff01101fa912409fa912509fe701109ffe01107ffc0012bfc50149cfff00101fef01001;
assign testcases[157] = 512'hfaa21697faa146a7fe702578fe901477fa915698f972678afff01001fff01101fa912409fa912509fe801109ffe01107ffc0012cfc50149cfff00101fef01001;
assign testcases[158] = 512'hfef00132fef00132ffe00123fff00122fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00016fff00125fff00001fff00000;
assign testcases[159] = 512'hfdf00233fdf01233ffd00223ffe00223fee01234fee11224fff00000fff00000fde00105fde00105ffe00004fff00003fff00016ffe00136fff00001fef00001;
assign testcases[160] = 512'hfef00122fef00122ffe00123fff00122fef01123fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00006fff00125fff00001fff00000;
assign testcases[161] = 512'hfdf10233fdf01233ffe00223ffe00223fee01234fee12224fff00000fff00000fde00105fde01105ffe00004fff00003fff00016ffe00136fff00001fef00001;
assign testcases[162] = 512'hfef00122fef00122ffe00123fff00122fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00016fff00125fff00001fff00000;
assign testcases[163] = 512'hfdf00233fdf01233ffe00223ffe00223fee01234fee11224fff00000fff00000fde00105fde01105ffe00004fff00003fff00016ffe00136fff00001fef00001;
assign testcases[164] = 512'hfef00132fef01132fff00122fff00122fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00015fff00125fff00001fef00001;
assign testcases[165] = 512'hfdf00133fdf01133ffe00233ffe00123fee01234fee01224fff00000fff00000fde00105fde00105ffe00004fff00003fff00016ffe00136fff00001fef00001;
assign testcases[166] = 512'hfef00122fef00122ffe00123fff00122fef01123fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00016fff00125fff00001fef00001;
assign testcases[167] = 512'hfdf00233fdf01233ffe00223ffe00223fee01233fee12224fff00000fff00000fde00105fde01205ffe00004fff00003fff00016ffe00126fff00001fef00001;
assign testcases[168] = 512'hfef00122fef00122fff00122fff00122fef01123fef01113fff00000fff00000fef00104fef00104fff00003fff00002fff00005fff00025fff00001fef00001;
assign testcases[169] = 512'hfdf00233fdf01233ffe00233ffe00123fee01233fee11224fff00000fff00000fde00105fde00105ffe00004fff00003fff00016ffe00136fff00001fef00001;
assign testcases[170] = 512'hfef00122fef00122ffe00123fff00122fef00123fef00123fff00000fff00000fef00004fef00104fff00003fff00003fff00016fff00025fff00001fef00001;
assign testcases[171] = 512'hfdf00233fdf01233ffd00233ffe00223fee01234fee11224fff00000fff00000fde00105fde01205ffe00004fff00003fff00016ffe00136fff00001fef00001;
assign testcases[172] = 512'hfef00043fef00043fff00033fff00033fef00044fff00034fff00000fff00000fef00005fef00004fff00004fff00003fff00016fff00046fff00001fff00001;
assign testcases[173] = 512'hfef00113fef00113ffe00134ffe00134fef00124fef00114fff00000fff00000fef00005fef00104ffe00005fff00004fff00007fff00016fff00001fef00001;
assign testcases[174] = 512'hfef00113fef01113ffc00235ffd00235fef01225fef11214fff00000fff00000fef00105fef00105ffc00006fff00005fff00007fff00116fff00001fef00001;
assign testcases[175] = 512'hfef00213fef01213ffb00346ffc00246fee12225fef12215fff00000fff00001fef00105fef00105ffb00107fff00106fff00007fff00116fff00001fef00001;
assign testcases[176] = 512'hfef00214fef01213ffa00347ffb00346fee01336fef12315fff00000fff00001fef00105fef00105ffa00108fff00107fff00007fff00116fff00001fef00001;
assign testcases[177] = 512'hfef10214fef01213fe901447fea01357fee12436fee12315fff00000fff00001fef00205fef00205ff900109ffe00107fff00007ffe00116fff00001fef00001;
assign testcases[178] = 512'hfef10314fef01214fe901447fea01457fee12436fee12415fff00000fff00001fef01205fef01205ff900109ffe00108fff00108ffe00116fff00001fef00001;
assign testcases[179] = 512'hfdf10324fdf12324fe801558fe901457fde23436fee23425fff00001fff00001fef01205fef01205fe80010affe00108fff00118ffe00217fff00001fef00001;
assign testcases[180] = 512'hfdf10324fdf02324fe701569fe801468fdd12447fee12426fef00001fff00001fdf01206fef01205fe70010bffe00109fff00118ffe00227fff00001fef00001;
assign testcases[181] = 512'hfdf11324fdf12324fe601669fe701569fdd13537fde13526fef00101fff01101fde11206fef01205fe60020cffd0010afff00118ffe00227fff00001fef00001;
assign testcases[182] = 512'hfde11424fde13424fe50177afe60167afdd14637fde14626fef01101fff01101fde11306fde01305fe40120dffd0020bfff00118ffe00227fff00101fef00001;
assign testcases[183] = 512'hfde21424fde13424fe40287bfe50177bfdd15747fdd24626fef01101fff01101fde11306fde11306fe30120effd0120cfff00119fed01327fff00101fef00001;
assign testcases[184] = 512'hfde11455fde13455fd4017bbfe5016cbfdd15797fdd24656fef01101fff01101fde11306fde11306fe30020effd0021cfff00129fed01358fff00101fef00001;
assign testcases[185] = 512'hfde21525fde13525fd30298bfd40189bfcc26847fdd25726fef11101fef11101fde11306fde11306fd20120effc0120cffe00119fed01328fff00101fef01101;
assign testcases[186] = 512'hfde21525fde14525fd202a9cfd30299cfcc26948fdd26726fef11101fef11101fde11406fde11406fd10130fffc0130cffe00119fec01328fff01101fef01101;
assign testcases[187] = 512'hfef00012fef00012fff00013fff00012fff00013fff00013fff00000fff00000fef00004fef00004fff00003fff00003fff00006fff00015fff00001fff00000;
assign testcases[188] = 512'hfef00113fef00113ffe00124ffe00123fef00124fef01114fff00000fff00000fef00104fef00104ffe00005fff00004fff00006fff00016fff00001fff00000;
assign testcases[189] = 512'hfef00113fef01113ffd00235ffd00134fef01225fef01214fff00000fff00000fef00105fef00104ffd00006fff00005fff00007fff00116fff00001fef00000;
assign testcases[190] = 512'hfef10223fef11223ffb01346ffb00246fee01335fef11325fff00000fff00000fef00105fef00105ffb00107fff00106fff00017fff00116fff00001fef00001;
assign testcases[191] = 512'hfef00223fef01223fea00356ffb00256fee02335fef11324fff00000fff00000fef00105fef00105ffa00108fff00106fff00017fff00116fff00001fef00001;
assign testcases[192] = 512'hfef10223fef01223fe901457fea01366fde12336fee12325fef00000fff00001fef00205fef00205fe900108ffe00107fff00017ffe00126fff00001fef00001;
assign testcases[193] = 512'hfef10224fef01223fe901457fea01367fee12436fee12425fff00000fff00001fef01205fef01205fe900109ffe00107fff00117ffe00126fff00001fef00001;
assign testcases[194] = 512'hfef00113fef01113ffc00235ffd00244fef01235fef01214fff00000fff00000fef00105fef00104ffc00106fff00005fff00007fff00116fff00001fef00000;
assign testcases[195] = 512'hfdf10324fdf12324fe801468fe901478fde12446fee12425fff00001fff00001fef01205fef01205fe80010affe00108fff00118ffe00227fff00001fef00001;
assign testcases[196] = 512'hfdf21324fdf12324fe701578fe801478fdd13546fee13425fef00001fff01101fdf11205fef01205fe70010bffe00109fff00118ffe00227fff00001fef00001;
assign testcases[197] = 512'hfde11424fde12324fe601679fe701589fdd14647fde14526fef01101fff01101fde11306fde01305fe50020cffd0020afff00118ffe00227fff00001fef00001;
assign testcases[198] = 512'hfde11424fde13424fe50178afe60168afdd15747fdd24626fef01101fff01101fde11306fde11305fe40120dffd0020bfff00118fed01227fff00101fef00001;
assign testcases[199] = 512'hfde11424fde13424fe40288bfe50179bfdc15747fdd25626fef01101fff01101fde11306fde11306fe30120effd0120bfff00119fed01328fff00101fef00001;
assign testcases[200] = 512'hfde21535fde15524fd30299bfd4028abfcc36857fdd46736fef11101fef11101fde11306fde11306fd20120effd0120cffe00119fed01328fff01101fef01101;
assign testcases[201] = 512'hfde21535fde14535fd20299cfd4029acfcc26958fdd26736fef11101fef11101fde11406fde12406fd20130fffc0120cffe00119fec01328fff01101fef01101;
assign testcases[202] = 512'hfef00012fef00012fff00012fff00012fef00013fef00013fff00000fff00000fef00004fef00004fff00003fff00003fff00006fff00015fff00001fff00000;
assign testcases[203] = 512'hfef00113fef00113ffe00123ffe00123fef00124fef01114fff00000fff00000fef00104fef00104ffe00004fff00004fff00006fff00016fff00001fff00000;
assign testcases[204] = 512'hfef00123fef01113ffc00245ffc00245fee01235fef01224fff00000fff00000fef00105fef00104ffc00107fff00106fff00017fff00116fff00001fef00001;
assign testcases[205] = 512'hfef00223fef01213ffb00346ffb00246fee01336fef12325fff00000fff00000fef00105fef00105ffb00108fff00106fff00017fff00116fff00001fef00001;
assign testcases[206] = 512'hfef10224fef01213fea01457ffa01357fee12336fef12325fff00000fff00001fef00205fef00205ffa00109ffe00107fff00017fff00116fff00001fef00001;
assign testcases[207] = 512'hfef10324fef01224fe901457fea01457fee12436fee12425fff00000fff00001fef01205fef01205fe900109ffe00108fff00118ffe00127fff00001fef00001;
assign testcases[208] = 512'hfdf11324fdf12324fe801558fe901468fde23436fee23425fff10000fff11001fef11205fef01205fe80010affe00108fff00118ffe00227fff00001fef00001;
assign testcases[209] = 512'hfdf11324fdf12324fe701568fe801468fdd13546fde13425fef00001fff00001fef01205fef01205fe60010bffe00109fff00118ffe00227fff00001fef00001;
assign testcases[210] = 512'hfdf11324fdf12324fe701669fe701579fdd13547fee13526fef00001fff01101fde11206fef01205fe60020cffd0010afff00118ffe00227fff00001fef00001;
assign testcases[211] = 512'hfde11424fde13424fe50177afe60168afdd14647fde14626fef01101fff01101fde11306fde01305fe40120dffd0020bfff00118fed00227fff00101fef00001;
assign testcases[212] = 512'hfde11424fde13424fe40187bfe50178bfdd15747fdd24626fef01101fff01101fde11306fde11306fe30120effd0120cfff00119fed01328fff00101fef00001;
assign testcases[213] = 512'hfde21525fde13424fd30298bfe40289bfdc15847fdd25726fef11101fff01101fde11306fde11306fe20120fffc0120cffe00119fed01328fff00101fef01101;
assign testcases[214] = 512'hfde11424fde13424fd30189bfd4017abfdd15757fdd24626fef11101fef01101fde11306fde11306fd20120fffc0120cffe00119fed01328fff00101fef01101;
assign testcases[215] = 512'hfde11424fde13424fe30188bfd40179bfcd15747fdd25626eef11101fef11101fde11306fde11305fd10120effc0120cffe00118fed01327fff00101fef01101;
assign testcases[216] = 512'hfef10113fef00113ffd00134ffd00134fef01125fef01114fff00000fff00000fef00104fef00104ffd00006fff00005fff00007fff00116fff00001fef00001;
assign testcases[217] = 512'hfef00012fef00012fff00013fff00012fef00013fff00013fff00000fff00000fef00004fef00004fff00003fff00003fff00006fff00015fff00001fff00000;
assign testcases[218] = 512'hfef00113fef00113ffe00124ffe00123fef00124fef00114fff00000fff00000fef00004fef00004ffe00005fff00004fff00006fff00015fff00001fff00000;
assign testcases[219] = 512'hfef00113fef00113ffd00234ffd00134fef01225fef01214fff00000fff00000fef00104fef00104ffd00006fff00005fff00007fff00116fff00001fef00001;
assign testcases[220] = 512'hfef00113fef01113ffc00245ffc00245fef01225fef01214fff00000fff00000fef00105fef00104ffc00107fff00106fff00007fff00116fff00001fef00001;
assign testcases[221] = 512'hfef00213fef01213ffb00346ffc00246fee01335fef11214fff00000fff00000fef00105fef00104ffb00107fff00106fff00007fff00116fff00001fef00001;
assign testcases[222] = 512'hfef10213fef01213ffa01356ffb00356fee12335fef12315fff00000fff00001fef00105fef00105ffa00108ffe00107fff00007fff00116fff00001fef00001;
assign testcases[223] = 512'hfef10223fef01213fea01457fea01357fee12436fef12325fff00000fff00001fef00205fef00205fe900109ffe00108fff00017ffe00116fff00001fef00001;
assign testcases[224] = 512'hfef10324fef02213fe901457fe901467fee12436fee12425fff00001fff00001fef01205fef01205fe80010affe00108fff00117ffe00116fff00001fef00001;
assign testcases[225] = 512'hfdf11324fdf12324fe801568fe801468fde23536fee13425fef10001fff11001fef11205fef01205fe70010bffe00109fff00118ffe00227fff00001fef00001;
assign testcases[226] = 512'hfdf10224fdf01224fe801478fe801378fde12446fee12425fef00001fff00001fdf01205fef01205fe70010bffe00109fff00118ffe00227fff00001fef00001;
assign testcases[227] = 512'hfdf11324fdf12324fe601679fe701579fdd14546fee13525fef01101fff01101fde11205fdf01205fe50020cffd0010afff00118ffe00227fff00101fef00001;
assign testcases[228] = 512'hfde11424fde13324fe50177afe60168afdd14647fde14525fef01101fff01101fde11306fde01305fe40120dffd0020bfff00118fee00227fff00101fef00001;
assign testcases[229] = 512'hfde11424fde13424fe40178afe50179bfdd16747fde25626fef01101fff01101fde11306fde11305fe20120effc0120cfff00118fed01327fff00101fef01101;
assign testcases[230] = 512'hfde21524fde13424fd30288bfd40179bfdd26847fdd25626fef11101fef01101fde11306fde11305fd20120fffc0120cfff00119fed01327fff00101fef01101;
assign testcases[231] = 512'hfde21524fde14524fd30299bfd40289cfcc26847fdd25726fef11101fef11101fde11306fde11306fd10130fffc0130dffe00119fed01328fff01101fef01101;
assign testcases[232] = 512'hfef00012fef00012fff00023fff00023fff00013fff00013fff00000fff00000fef00004fef00004fff00004fff00003fff00006fff00015fff00001fff00000;
assign testcases[233] = 512'hfef00113fef00113ffe00124ffe00123fef00124fef00114fff00000fff00000fef00004fef00004ffe00005fff00004fff00006fff00015fff00001fff00000;
assign testcases[234] = 512'hfef00113fef00113ffd00235ffd00134fef01225fef01114fff00000fff00000fef00104fef00104ffd00006fff00005fff00006fff00116fff00001fef00001;
assign testcases[235] = 512'hfef00113fef01113ffc00235ffc00245fef01225fef01214fff00000fff00000fef00105fef00104ffc00107fff00106fff00007fff00116fff00001fef00001;
assign testcases[236] = 512'hfef10213fef01213ffb01346ffb01346fee02325fef11214fff00000fff00000fef00105fef00104ffb00108fff00107fff00007fff00116fff00001fef00001;
assign testcases[237] = 512'hfef10213fef01213ffa01447ffb01346fee12335fef12315fff00000fff00001fef00105fef00105ffa00108ffe00107fff00007fff00116fff00001fef00001;
assign testcases[238] = 512'hfef10213fef01213fe901457fea01357fde12436fef12315fff00000fff00001fef00205fef00205fe900109ffe00108fff00007fff00116fff00001fef00001;
assign testcases[239] = 512'hfef11324fef02214fe801558fe901458fde13436fee22425fef10001fff01001fef11205fef01205fe70010affe00109fff00118ffe00116fff00001fef00001;
assign testcases[240] = 512'hfdf11324fdf12324fe801568fe801468fee13536fee13425fff00001fff00001fef01205fef01205fe70010bffe00109fff00118ffe00217fff00001fef00001;
assign testcases[241] = 512'hfdf11324fdf12324fe701669fe701569fde13536fee13425fef00001fff01101fef01205fef01205fe60020cffd0010afff00118ffe00227fff00001fef00001;
assign testcases[242] = 512'hfdf11424fdf12324fe60166afe60167afdd14637fde14525fef01101fff01101fde11205fdf01205fe40020dffd0020bfff00118ffe00227fff00101fef00001;
assign testcases[243] = 512'hfde11424fde13424fe40177afe50178bfdd15747fde24626fef01101fff01101fde11306fde11305fe20120effc0120cfff00118fed01227fff00101fef00001;
assign testcases[244] = 512'hfde11424fde13424fe40287bfd40178bfdd15747fdd25626fef01101fff01101fde11306fde11305fd10120fffc0120dfff00119fed01327fff00101fef01101;
assign testcases[245] = 512'hfde21524fde14424fd20298cfd30289cfdc26847fdd25726fef11101fef11101fde11306fde11306fd00130fffc0120dffe00119fed01328fff00101fef01101;
assign testcases[246] = 512'hfde21525fde14524fd202a8cfd30299cfcc27948fdd26726fef11101fef11101fde11406fde11306fd00130fffc0130effe00119fed01328fff01101fef01101;
assign testcases[247] = 512'hfde00001fde00001fd200102fd300101fdc00002fdd00002fef00000fef00000fde00003fde00003fd000002ffc00002ffe00004fed00004fff00001fef00000;
assign testcases[248] = 512'hfde11323fde12323ffb01556ffb01556fee12334fee12324fdd23313fed13313fde11205fde01205ffb00106fff00105fff00016ffe00126fed01303fde02203;
assign testcases[249] = 512'hfcd11344fcd13344fe702678fe802578fdd12345fdd13335ecb35525fdc24424fcc11306fcc11306fe801109ffe01108ffe00017fec00247fec02405fcc14404;
assign testcases[250] = 512'hfef10223fef01123ffc01334ffd01344fef01123fef01223fee12212fee12212fef00104fef01104ffd00105fff00104fff00015fff00125ffe01202fee02202;
assign testcases[251] = 512'hfcd22656fcd25556fea1498afeb1389afdd35557fdd45547eef67726fef46625fcd42408fcd32408ffb0120bffe0120afff00119fec01248fff14605eef26505;
assign testcases[252] = 512'heab21657eab24657fe61398afe71389afbb14557ebb24547db947726eca36625ebb12408dab12508fe60120bffd0120affe00119eda01259edb14605ebb16505;
assign testcases[253] = 512'hfde11213fde12213ffd01323ffe01223fee12213fee12313fff00000fff00000fde11204fde01204ffd00104fff00103fff00006ffe00115fff00001fef00000;
assign testcases[254] = 512'hfbb32857fbb27767fe802868fe902677fb927869fb938968fff00001fff01101fba23609fba23709fe901209ffe01208ffc0112bfd70156bfff00101fef00001;
assign testcases[255] = 512'hfcc32756fcc27766fea02667fea02677fba26767fba37858fff00001fff00101fcb23608fcb23608ffa01208ffe01207ffd0112afd90146afff00101fef00001;
assign testcases[256] = 512'hfbc32766fbc27766fea02767fea02667fba26777fba37858fff00001fff00101fbb23608fbb13608fe901208ffe01207ffd0112afd90146afff00101fef00001;
assign testcases[257] = 512'hfde10223fde02223ffd01234ffe01233fee02224fee12324fff00000fff00000fde01205fde01205ffe00104fff00104fff00016ffe00126fff00001fef00001;
assign testcases[258] = 512'hfbb32756fbb27766fe902667fea02667fba26768fba37858fff00001fff00101fba23508fbb13608fe901208ffe01207ffd0112afd80146afff00101fef00001;
assign testcases[259] = 512'hfde10223fde01223ffd01234ffe01233fee02234fee12324fff00000fff00000fde01205fde01205ffd00104fff00104fff00016ffe00136fff00001fef00001;
assign testcases[260] = 512'heab32756fab26756fe802667fe902677ea926768da937858fff00001fff00001eaa23508daa13608fe901208ffe01207ffd0012afc80146afff00101fef00001;
assign testcases[261] = 512'hfab32736fab26736fe702857fe812857fba15636faa26726fff12201fff13201faa22507faa12608fe801208ffe01207ffd00119fd901338fff02201fef12201;
assign testcases[262] = 512'hfbb32646fbb26646fe802667fe902667fba26747fba37737fff00000fff00001fba23508fba13608fe801208ffe01207ffd0011afd801449fff00101fef00001;
assign testcases[263] = 512'hfbb32746fbb26646fe802667fe902677fba26757fba37847fff00000fff00001fba23508fba13608fe801208ffe01207ffd0011afd80144afff00001fef00001;
assign testcases[264] = 512'hfce32814fce26813fe502c7afe602b7afdd27b26fdd37a15fee58701fee49701fcd22706fde13705fe50130cffd0130affe01218fed01527fee16801fef27601;
assign testcases[265] = 512'hfde11414fce13413fd302a8bfd40299bfdd15726fdd24615fee12201fee12201fde12406fde12405fd20130dffc0130cffe00118fed01327ffe01202fef01101;
assign testcases[266] = 512'hfde11414fde13413fd20298bfd30299bfcd15726fdd24615eee12201fee12201fde12406fde12405fd10130effc0120cffe00118fed01327fef01101fef01101;
assign testcases[267] = 512'hfde11424fce13424fd30298cfd30289cfdd15736fdd24525fee11111fee11101fdd11306fde11306fd20130effc0130cffe00119fed01327ffe01102fef01101;
assign testcases[268] = 512'hfde11424fde13424fd30298bfd40289cfdd15736fdd24525fef11201fef11101fde11406fde11305fd20130effc0120cffe00118fed01327fff01101fef01101;
assign testcases[269] = 512'hfde21424fde13414fd212b8cfd302a9cfcc68736fdd66625fee32211fee32211fdd42406fde32406fd11130effc1130cffe01119fec01327fee11102fef11101;
assign testcases[270] = 512'hfde11424fde14424fd30298cfd30299cfdd25736fdd34525fee21101fee12101fde12406fde21306fd20130effc0130cffe00119fed01327fff01101fef01101;
assign testcases[271] = 512'hfef00012fef00012fff00122fff00122fff00012fff00012fef11112fee01112fef00003fef00003fff00003fff00002fff00005fff00014ffe01102fef01102;
assign testcases[272] = 512'hfef00112fef00112ffe00123fff00122fef00112fef00112fdd12213fed12213fef00004fef00104fff00003fff00003fff00005fff00015fed01203ede01203;
assign testcases[273] = 512'hfef00122fef01122ffe00223ffe00233fef01123fef01113edd23313fdd13314fef00104fef00104ffe00004fff00003fff00005fff00025fed02304fdd12203;
assign testcases[274] = 512'hfef00122fef01122ffe00233ffe00233fef01123fef01113ecc24414fdc24414fef00104fef00104ffe00004fff00003fff00005fff00025fec02404fcd13304;
assign testcases[275] = 512'hfef00123fef01122ffd01334ffe01233fef01123fef01123ecb24414fdb24415fef00104fef00104ffe00104fff00104fff00015fff00125fdb03405fcc14404;
assign testcases[276] = 512'hfdf10233fdf01133ffc01344ffd01344fef01133fef01223eba36625fca36615fde00105fde00105ffd00105fff00104fff00016ffe00125fda13606ebb15505;
assign testcases[277] = 512'hfde10233fde01233ffc01345ffd01344fee01234fee11234ea947726fc937726fde00105fde01205ffc00105fff00105fff00016ffe00136fc914607eba16606;
assign testcases[278] = 512'hfde10244fde01243ffb01455ffc01355fde01244fde12234ea948827eb838827fde01205fde01205ffc00106fff00105fff00016fed00136ec815707eaa27706;
assign testcases[279] = 512'hfce10244fde02244feb01456ffc01455fde01244fdd12234e9858828eb848828fdd01206fdd01206ffb00106fff00105fff00017fed00146ec815808ea927707;
assign testcases[280] = 512'hfcd10254fcd02254fea01466feb01366fdd02244fdd12245e9759828ea749828fcd01206fcd01206ffb00107fff00106fff00017fed00147ec716808ea928707;
assign testcases[281] = 512'hfcd11354fcd12354fea01466fea01466fdd02345fdd12345d9759928ea74a929fcd11206fcc01206fea01107ffe00106ffe00017fec00147eb716909e9828808;
assign testcases[282] = 512'hfcd11355fcc12355fe901567fea01476fcc02355fcc12345d875aa29ea64aa29fcc11206fcc01306fe901108ffe00107ffe00017fec00257eb616a09d9829908;
assign testcases[283] = 512'hfbc11355fbc12365fe801577fe901477fcc12355fcc12345d866aa29ea65ba29fcc11207fbc01307fe901108ffe00107ffe00018feb00257eb617a0ad972a909;
assign testcases[284] = 512'hfbc11365fbc12365fe801477fe901477fcb12365fcb12356c767ca2ad966ca2afbb11207fbb01307fe801108ffe01107ffe00018feb00258da617a0ad873b909;
assign testcases[285] = 512'hfab11466fab12466fe701578fe801488fbb12366fbb12456d867ca2ae955cb2afbb11307fba01308fe701109ffe01108ffe00018fda00268eb618b0ad873ba09;
assign testcases[286] = 512'hffb11466ffb12366ff701578ff801478ffb12366ffb12356ff67cb2aff56cb2affb11308ffa01308ff701109ffe01108ffe00018ffa00268ff618b0aff73ba09;
assign testcases[287] = 512'hfab11465fab12466fe701578fe801477fbb12366fbb12456c866aa2ad965ba2afab11307fab01307fe801109ffe01108ffe00018fda00258db617a0ad972a909;
assign testcases[288] = 512'hfbc11455fbc12365fe801577fe901477fcc12355fcc12346d876aa29ea65ba29fbb11307fbb01307fe801108ffe00107ffe00018feb00258eb617a09d9829909;
assign testcases[289] = 512'hfef00012fef00012fff00112fff00112fff00012fff00012fee11102fee01102fef00003fef00003fff00003fff00002fff00005fff00014ffe01102fef01102;
assign testcases[290] = 512'hfef00112fef00012ffe00123fff00123fef00112fef00112edd12213fed12213fef00004fef00004fff00003fff00003fff00005fff00015fed01203ede02202;
assign testcases[291] = 512'hfef00122fef00122ffe00223ffe00223fef00113fef01113edd23313edd13314fef00104fef00104ffe00004fff00003fff00005fff00025fed02304edd12203;
assign testcases[292] = 512'hfef00122fef01122ffd00234ffe00233fef01123fef01123ecc24414fdc24414fef00104fef00104ffe00104fff00103fff00015fff00025edc02404ecd13304;
assign testcases[293] = 512'hfef00123fef01123ffd01334ffe01234fef01123fef01123ecc24414fdb24415fef00104fef00104ffd00104fff00104fff00015fff00125fdb03405ecc14404;
assign testcases[294] = 512'hfde00233fdf01233ffc01344ffd01344fee01233fee01223daa36515fba36615fde00105fde00105ffd00105fff00104fff00016ffe00136fca13606ebb15505;
assign testcases[295] = 512'hfde10233fde01233ffc01445ffc01345fee01234fee11234eba47626ec937716fde00205fde01205ffc00106fff00105fff00016ffe00136ec914707eba16506;
assign testcases[296] = 512'hfde10244fde01244ffb01455ffc01355fde01244fde11234d9947727eb837727fde01205fdd01205ffb00106fff00105fff00016fed00136ec914707eaa26606;
assign testcases[297] = 512'hfcd10344fcd02344fea01456ffb01456fdd01244fdd12335d9858827da848828fcd01206fcd01206ffb00107fff00106fff00017fed00147eb815808d9927707;
assign testcases[298] = 512'hfcd11344fcd12354fea01556fea01466fdd02345fdd12345e9859928eb749928fcd01206fcc01306fea00107ffe00106ffe00017fec00147ec815908ea928807;
assign testcases[299] = 512'hfcd11355fcd12355fe901567fea01466fdd02355fcc12345c7759928d9649929fcc01206fcc01306fea00108ffe00106ffe00017fec00247eb616909d9828808;
assign testcases[300] = 512'hfbc11355fbc12355fe901567fea01467fcc02355fcc12345c7759a29d9649a29fcc11307fbc01307fe901108ffe01107ffe00018feb00257db616a09d8828908;
assign testcases[301] = 512'hfef00012fef00012fff00012fff00012fff00012fff00012fee11103fee01103fef00003fef00003fff00003fff00002fff00005fff00014fee00103fef01103;
assign testcases[302] = 512'hfef00012fef00012fff00123fff00023fff00013fef00012edd21215fdc21205fef00004fef00004fff00003fff00003fff00005fff00015fec01205edd01104;
assign testcases[303] = 512'hfef00012fef00012ffe00123ffe00123fef00013fef00013ecb22316fcb12316fef00004fef00004ffe00004fff00003fff00005fff00015fdb01306ecc12205;
assign testcases[304] = 512'hfef00123fef00123ffe00134ffe00134fef00123fef00113eba23417eca23417fef00004fef00104ffe00004fff00004fff00005fff00025eda02408ebb13307;
assign testcases[305] = 512'hfdf00123fdf00123ffd00234ffe00134fef00123fef11123ea975518eb925518fef00105fef00105ffd00005fff00004fff00016ffe00025ec903509eaa34508;
assign testcases[306] = 512'hfde00123fde00123ffd00234ffd00244fee01124fee01124d9835619eb735619fde00105fde00105ffd00005fff00004fff00016ffe00026ec813609ea915608;
assign testcases[307] = 512'hfde00124fde01124ffc00235ffd00245fde01124fde01124c8736619da73661afde00105fde00105ffd00006fff00005fff00016fee00126eb71360ac9815609;
assign testcases[308] = 512'hfde00124fde01124ffc00245ffd00245fee01134fee01124d874771ae973671afde00105fde00105ffc00106fff00105fff00016ffe00136eb71470ad8826709;
assign testcases[309] = 512'hfcd00234fdd01234ffb00346ffc00345fdd01235fdd01235d865891bea54891bfdd00106fdd00206ffc00106fff00106fff00017fed00137eb61590bd872780a;
assign testcases[310] = 512'hfcc10235fcc01245ffa01356ffb01356fdc01245fdc11236d7459a1cd8449a1cfcc00207fcc01207ffb00107fff00106ffe00018fec00148da415a0cc752990b;
assign testcases[311] = 512'hfbc10346fcc01345fea01457fea01357fcc01346fcc12336b546bb1dc735bb1dfcc01207fcb01307ffa00108ffe00107ffe00018feb00148d9316b0dc553ab0c;
assign testcases[312] = 512'hfab10457fab12457fe801468fe901468fbb12357fbb12447a527cc2ec726cc1efba01308faa01308fe900109ffe00108ffe00019fda00259d9217c0eb433bc0e;
assign testcases[313] = 512'hfaa11557faa12567fe801568fe801478fba12467fba12457a418ee2fc717ee1ffba11309fa901409fe800109ffe00108ffd00119fd900259d9118e0fa424ee0f;
assign testcases[314] = 512'hf9911568fa913568fe701579fe801589fb912568fb9135589209ff2fb507ff1ffa911409fa91140afe70010affe00108ffd0012afd80026ac8029f0f9314ff0f;
assign testcases[315] = 512'hfef00012fef00012fff00012fff00012fff00012fff00012fef00013fee00003fef00003fef00003fff00003fff00002fff00005fff00014ffe00003fef00003;
assign testcases[316] = 512'hfef00012fef00012fff00123fff00023fef00013fef00013edd11115fdc11215fef00004fef00004fff00004fff00003fff00005fff00015fec01205edd01104;
assign testcases[317] = 512'hfef00013fef00012ffe00123ffe00123fef00013fef00013ecb12316edb12316fef00004fef00004ffe00004fff00003fff00005fff00015fdb01306ecc12205;
assign testcases[318] = 512'hfef00123fef00123ffe00134ffe00134fef00123fef00113eba23417eca23417fef00005fef00105ffe00005fff00004fff00006fff00025eda02408ebb13307;
assign testcases[319] = 512'hfde00123fdf00123ffd00234ffd00134fee00124fee00124ea934518eb834518fde00105fde00105ffd00005fff00004fff00016ffe00026ec912509eaa14408;
assign testcases[320] = 512'hfde00124fde01124ffc00235ffd00235fee01124fde01124d9835619eb725619fde00105fde00105ffd00006fff00005fff00016ffe00126ec71360ada915509;
assign testcases[321] = 512'hfde00124fde01124ffc00235ffc00245fde01134fde01124d874671aea73671afde00106fdd00106ffc00106fff00105fff00017fed00136eb71470ad9826609;
assign testcases[322] = 512'hfcd00234fdd01234ffb00346ffc00245fdd01235fdd01225d864781ada63781bfdd00106fdd00106ffc00106fff00105fff00017fed00137eb61480bd872770a;
assign testcases[323] = 512'hfcd00235fcd01235ffb01346ffb01346fdd01235fcd01235c755991bd9549a1bfcd00206fcc00207ffb00107fff00106fff00017fec00137da515a0cc762890b;
assign testcases[324] = 512'hfcd10335fcd01335ffb01446ffb01356fdd01235fdc11335d756aa1cd945ab1cfcc01207fcc01207ffb00107fff00106ffe00017fec00137ea516b0cd7639a0b;
assign testcases[325] = 512'hfbb10346fbb12346fe901457fea01457fcb02346fcb12336b637bc1dd835bc1dfcb01208fbb01308ffa00108ffe00107ffe00018feb00248da316c0dc643bb0d;
assign testcases[326] = 512'hfaa11457faa12457fe801468fe901468fba02357fba12447a527cc2fc726cd1ffaa01308faa01309fe800109ffe00108ffd00019fd900259c9217d0fb423cc0e;
assign testcases[327] = 512'hfa911558fa913558fe701568fe801578fa912558fa9135489419ff1fc717ef1ffa911409fa911409fe80010affe00108ffd0011afd80025ac9128f0fb414ff0f;
assign testcases[328] = 512'hf9911658f9913668fe601579fe701579e9813568f9813658900aff1fc407ff1ff981140af981150afe60010affd00109ffc0011aec70036ac6029f0fa004ff0f;
assign testcases[329] = 512'hfef00012fef00012fff00012fff00012fff00012fff00012eee11103fee01103fef00003fef00003fff00003fff00002fff00005fff00014ffe00103fef01103;
assign testcases[330] = 512'hfef00012fef00012fff00123fff00123fef00013fef00013edc32215fdc22205fef00004fef00004fff00004fff00003fff00005fff00015fec11205edd02204;
assign testcases[331] = 512'hfef00113fef00113ffe00124ffe00123fef00113fef00113dbb22316ecb12316fef00004fef00004ffe00004fff00004fff00005fff00015edb01306ebc12305;
assign testcases[332] = 512'hfdf00113fdf00123ffd00124ffe00134fef00123fef00113eba24417ec924417fef00105fee00105ffe00005fff00004fff00006ffe00026ec902408ebb13407;
assign testcases[333] = 512'hfde00124fde00124ffd00235ffd00235fee01124fee01124da934518eb824518fde00105fde00105ffd00005fff00005fff00016ffe00126ec803508eaa14507;
assign testcases[334] = 512'hfde00224fde01124ffc00235ffc00235fde01124fde01224d9835619eb735619fde00106fdd00106ffc00106fff00105fff00017fed00126ec813609da915608;
assign testcases[335] = 512'hfdd00224fdd01224ffc00335ffc00245fdd01225fdd01225d974671aea73671afdd00106fdd00206ffc00106fff00105fff00017fed00127eb71470ad9826709;
assign testcases[336] = 512'hfcd00235fcd01235ffb00346ffc00246fdd01235fdd01225d864671aea63671bfdd00106fdd00106ffc00107fff00106fff00017fed00137eb61470bd872670a;
assign testcases[337] = 512'hfcc10335fcc01335ffa01446ffb01346fdc01236fdc11336c755891bd954891cfcc00207fcc01207ffb00107fff00106ffe00018fec00138da51590cc762890b;
assign testcases[338] = 512'hfbb10336fbb12346fe901447fea01457fcb12346fcb12336b646ab1dd835ab1dfbb01308fbb01308fe900108ffe00107ffe00018fea00239d9316b0dc643aa0c;
assign testcases[339] = 512'hfbb11436fbb12446fe901557fea01457fcb12446fcb12437c637cc1dd836cc1dfbb11308fbb01408fe900108ffe00107ffe00119fda00239d9317c0dc543bc0c;
assign testcases[340] = 512'hfaa11447faa12458fe801558fe901468fba12458fba12448b427cd1ec726dd1efaa11309fa901409fe80010affe00108ffd0011afd90024ad9217d0fa523cd0e;
assign testcases[341] = 512'hf9911658f9913658fe701669fe801579fa913558fa913649a419ee1fc717ef1ffa91140af981150afe70010affe00109ffd0011afd80035bc8128f0f9314ee0f;
assign testcases[342] = 512'hd8811759d8813769fe60167afe70157afa813669ea813659930aff1fb607ff1fe981150bd971260bfe60020bffd00209ffc0011bfc60136bb8029f0fa304ff0f;
assign testcases[343] = 512'hf8811759f9813769fe60167afe70157afa713669fa8136599309ff1fb607ff1ff971150bf971260bfe60020bffd00109ffc0011bfc60136bc8029f0f9314ff0f;
assign testcases[344] = 512'hf9921658f9913669fe701579fe801579fa813559fa923659a319fe1fb61afe1ffa81140af981150afe70010affe00109ffd0011afd70035bc8128f0fa416fe0f;
assign testcases[345] = 512'hfaa10368faa01378fe801478fe801379fb902378fba12358b5269a2fc7249a2ffa901209fa90130afe80010affe00108ffd0002afd90026ad9216a0fb5229a0f;
assign testcases[346] = 512'heaa10377eba01387fe800378fe900278fba01277fba11367b633673ec823673ffba00209fba01209fe900109ffe00108ffd00029fd900179d931370fb532670e;
assign testcases[347] = 512'hfbb10346fbb12347fe901457fea01457fbb02347fbb12337b646aa1dd835ab1dfbb01308fba01308fe900108ffe00107ffe00019fda00249da416b0dc643aa0c;
assign testcases[348] = 512'hfcc10336fcc01336ffa01447ffb01347fcc01336fcc11336c755991bd844991cfcc01207fcc01207ffa00108fff00107ffe00018feb00138ea51590cd762890b;
assign testcases[349] = 512'hfcd00235fcd01235ffb00346ffc00346fdd01235fdd01225d864781ada63781afcd00207fcc00207ffb00107fff00106ffe00017fec00137eb61480bd972770a;
assign testcases[350] = 512'hfcd00225fdd01225ffb00336ffc00246fdd01225fdd01225d8746719da736719fdd00106fdd00206ffc00107fff00106fff00017fed00127eb71470ad9816609;
assign testcases[351] = 512'hfde00224fde01224ffc00235ffc00235fde01125fde01225d9835619eb835619fdd00106fdd00106ffc00106fff00105fff00017fed00127ec813609ea915508;
assign testcases[352] = 512'hfde00124fde01124ffc00235ffd00235fee01124fee01124ea934518eb824518fde00106fde00106ffd00006fff00005fff00016ffe00126ec902508eaa14507;
assign testcases[353] = 512'hfde00113fdf00123ffd00224ffd00134fee00124fee01114eba23417eca23417fde00105fde00105ffd00005fff00004fff00006ffe00026eda02407ebb13406;
assign testcases[354] = 512'hfdf00113fdf00113ffe00124ffe00124fef00113fef00113ecb22316ecb12316fef00105fdf00105ffe00005fff00004fff00006fff00016edb01306ecc12305;
assign testcases[355] = 512'hfef00013fef00012ffe00123fff00123fef00013fef00013ecd12204fdc12205fef00004fef00004fff00004fff00003fff00005fff00015edc01205ecd01204;
assign testcases[356] = 512'hfef00012fef00012fff00012fff00012fff00012fff00012fee11103fee01103fef00004fef00004fff00003fff00003fff00005fff00014ffe00103fef01103;
assign testcases[357] = 512'hfef00012fef00012fff00012fff00012fff00012fff00012fee11103fee01103fef00004fef00004fff00003fff00003fff00005fff00015fee00103fef01103;
assign testcases[358] = 512'hfef00013fef00012ffe00123fff00123fef00013fef00013edd11215fdc11215fef00004fef00004fff00004fff00003fff00005fff00015fec01205edd01104;
assign testcases[359] = 512'hfef00113fef00113ffe00124ffe00124fef00113fef00113ecb12316ecb12316fef00005fef00005ffe00005fff00004fff00006fff00015edb01306ecc12206;
assign testcases[360] = 512'hfde00123fdf00123ffd00224ffd00134fee00124fee00114daa23417eb923417fde00105fde00105ffd00005fff00004fff00006ffe00026ec902408ebb13407;
assign testcases[361] = 512'hfde00124fde01124ffc00235ffd00235fee01124fee01124da934518eb824518fde00106fde00106ffd00106fff00005fff00017ffe00126ec803509ea914508;
assign testcases[362] = 512'hfde00224fde01224ffc00335ffc00235fdd01225fdd01225c8835619da735619fdd00106fdd00106ffc00106fff00105fff00017fed00127eb713609d9815608;
assign testcases[363] = 512'hfcd00225fcd01225ffb00336ffc00336fdd01235fdd01225d874671aea63671afdd00206fdd00207ffc00107fff00106fff00017fed00137eb71470ad9826709;
assign testcases[364] = 512'hfcd10235fcd01235ffb01346ffb01346fdd01235fdd11225d864781ada63781bfcc00207fcc01207ffb00107fff00106ffe00018fec00138eb61480bd872780a;
assign testcases[365] = 512'hfbc10336fcc02336ffa01447ffb01447fcc02336fcc12336c7559a1bd9549a1cfcc01207fcb01308ffa00108ffe00107ffe00018feb00238ea515a0cc762990b;
assign testcases[366] = 512'hfbb11436fbb12446fe901547fea01457fcb12347fcb12437c546ab1cd745ab1cfbb01308fbb01308fea00108ffe00107ffe00019fea00249d9416b0cc653ab0c;
assign testcases[367] = 512'hfaa31547faa22447fe811558fe901558fba12447fba22438b63dcc1dc83ccc1efba11309fa911409fe900109ffe00108ffd0011afd90024ad9337c0eb636cc0d;
assign testcases[368] = 512'hf9911548fa913558fe701669fe801569fb913558fa913548b428dd1ec726dd1efa91140afa81150afe80010affe00109ffd0011afd80035ad9218d0fa523dd0e;
assign testcases[369] = 512'hd8811659d8813659fe601669fe701579e8813659d8813649a218ee1fb517ef1fe871150bd871150bfe60020bffd00109ffc0011beb60135bb7128f0f9214ee0f;
assign testcases[370] = 512'hf872175ae871476afe60167afe60167af971476af971475aa409ff1fc607ff1ff971150be861260cfe60020bffd0020affc0011cfc60136cc8029f0f8314ff0f;
assign testcases[371] = 512'hfdf00133fef01133ffd00244ffd00244fef01133fef01123fdd23314fed24414fef00104fef00104ffd00104fff00104fff00015fff00025fed02304fde13303;
assign testcases[372] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef01112ecd24414fdc24415fef00104fef00104ffe00104fff00003fff00005fff00015fec02405edd13304;
assign testcases[373] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef00112edd24414fdc25515fef00104fef00104ffe00004fff00003fff00005fff00025fec03405fdd14304;
assign testcases[374] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef00113ecc24525edc25515fef00104fef00104ffe00004fff00003fff00005fff00025edc03505edd14404;
assign testcases[375] = 512'hfef00122fef00122ffd00234ffe00233fef01123fef01113edc35525fdb25515fef00104fef00104ffe00104fff00003fff00005fff00025fec03505edd14404;
assign testcases[376] = 512'hfef00123fef00122ffd00234ffe01233fef01123fef01113edc35525edb25526fef00104fef00104ffe00104fff00103fff00005fff00025edc13505edd14404;
assign testcases[377] = 512'hfdf00123fef00122ffd00234ffd01244fef01123fef01113edc35525edb25526fef00104fef00104ffe00104fff00004fff00005fff00025edc13505edd14404;
assign testcases[378] = 512'hfef00123fef01122ffd00234ffd01244fef01123fef01123edc35525fdb25526fef00104fef00104ffe00104fff00104fff00015fff00025fec13506fdd14404;
assign testcases[379] = 512'hfdf00123fdf01122ffd01344ffd01244fee01123fef01123ecc36525ecb36626fdf00104fdf00104ffd00104fff00104fff00015fff00025edc13606ecd15404;
assign testcases[380] = 512'hfef00012fef00012fff00122fff00122fff00012fff00012eee12212fee12213fef00003fef00003fff00003fff00002fff00004fff00014fee01203fef01102;
assign testcases[381] = 512'hfef00112fef00012ffe00223fff00233fff00112fff00112edd23314fdd23314fef00004fef00004fff00003fff00003fff00005fff00014fed02304ede13303;
assign testcases[382] = 512'hfef00122fef00112ffe00233ffe00233fef00123fff00112edd24414fdc24414fef00004fef00104ffe00004fff00003fff00005fff00014fed02404fde13303;
assign testcases[383] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef00112edd24414edc24415fef00104fef00104ffe00004fff00003fff00005fff00015fec02405edd13304;
assign testcases[384] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef00113edd24414fdc25515fef00104fef00104ffe00004fff00003fff00005fff00025fec03405edd14304;
assign testcases[385] = 512'hfef00122fef01122ffe00233ffe01233fef01123fef01113edc35524fdc25525fef00104fef00104ffe00104fff00003fff00005fff00025fec03505edd14404;
assign testcases[386] = 512'hfef00123fef01122ffe01234ffe01233fef01123fef01113edc35525fdb25525fef00104fef00104ffe00104fff00103fff00005fff00025fec13505fdd14404;
assign testcases[387] = 512'hfdf00123fdf01122ffd01334ffd01234fef01123fef01113ecc35525edb26526fdf00104fdf00104ffd00104fff00103fff00005fff00025edc13505edd14404;
assign testcases[388] = 512'hfdf00123fef01122ffd01334ffd01234fef01123fef01113edc35525fdb36626fef00104fef00104ffe00104fff00104fff00015fff00025edc13505edd14404;
assign testcases[389] = 512'hfdf00123fef01122ffd01334ffd01234fef01123fef01123edc35525edb36626fef00104fef00104ffe00104fff00104fff00015fff00125eec13506edd15404;
assign testcases[390] = 512'hfdf10123fdf01122ffd01334ffd01244fef11123fef11123edca7625edb37626fef00104fef10104ffe00104fff00104fff00015fff00125eec14606edd46504;
assign testcases[391] = 512'hfef00123fef01122ffd01334ffd01244fef01123fef01123ecc36625fdb36626fef00104fef00104ffd00104fff00104fff00015fff00125fec14606fdd15505;
assign testcases[392] = 512'hfef00001fef00001fff00112fff00012fff00002fff00002fef01101fff01102fef00003fef00003fff00002fff00002fff00004fff00014fff00102fef01101;
assign testcases[393] = 512'hfef00012fef00012fff00122fff00122fff00012fff00012fee12212fee12213fef00003fef00003fff00003fff00002fff00004fff00014ffe01203fef01102;
assign testcases[394] = 512'hfef00012fef00012fff00122fff00122fff00012fff00012ede12213fed12313fef00003fef00003fff00003fff00002fff00005fff00014fee01203ede02202;
assign testcases[395] = 512'hfef00012fef00012fff00123fff00122fff00012fff00012edd23313fdd13314fef00003fef00003fff00003fff00003fff00005fff00014fed02304fde12203;
assign testcases[396] = 512'hfef00112fef00012fff00223fff00123fff00112fff00012edd23314fdc24414fef00003fef00003fff00003fff00003fff00005fff00014fed02304ede13303;
assign testcases[397] = 512'hfef00122fef00112ffe00223ffe00233fef00122fef00112edd24414fdc24414fef00004fef00104fff00003fff00003fff00005fff00014eed02404ede13303;
assign testcases[398] = 512'hfef00122fef00122ffe00233ffe00233fef00123fef00112edd24414edc24415fef00104fef00104ffe00004fff00003fff00005fff00015fec03405edd13304;
assign testcases[399] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef01113edd24414fdc25515fef00104fef00104ffe00004fff00003fff00005fff00025fec03405edd14404;
assign testcases[400] = 512'hfef00122fef01122ffe00233ffe00233fef01123fef01113ecc35515edc25515fef00104fef00104ffe00104fff00003fff00005fff00025edc03505ecd14404;
assign testcases[401] = 512'hfef00123fef01122ffe01234ffe01233fef01123fef01113ecc35525ecb25515fef00104fef00104ffe00104fff00103fff00005fff00025edc13505ecd14404;
assign testcases[402] = 512'hfef00123fef01122ffd00234ffe01234fef01123fef01113ecc35525edb25526fef00104fef00104ffe00104fff00103fff00005fff00025edc13505ecd14404;
assign testcases[403] = 512'hfef00133fef01132ffd01334ffe01244fef01133fef01123ecc35535edb25536fef00104fef00104ffe00104fff00104fff00015fff00025eec13506edd14404;
assign testcases[404] = 512'hfdf00123fef01122ffd01334ffd01234fef01123fef01123ecc35525edb25626fef00104fef00104ffe00104fff00104fff00015fff00125edc13506ecd14404;
assign testcases[405] = 512'hfdf00123fdf01122ffd01234ffd01244fef01123fef01123edc35525edb25626fdf00104fdf00104ffd00104fff00104fff00015fff00025eec13506edd15405;
assign testcases[406] = 512'hfdf00123fdf01122ffd01334ffd01244fee01133fef01123ecc35525edb36626fdf00104fdf00104ffd00104fff00104fff00015fff00125edc13606ecd15505;
assign testcases[407] = 512'hfef00012fef00011fff00012fff00012fff00012fff00012fef01112fff01112fef00003fef00003fff00003fff00002fff00004fff00014fff00102fef00102;
assign testcases[408] = 512'hfef00012fef00012fff00122fff00122fff00012fff00012eee12212fee12212fef00003fef00003fff00003fff00002fff00005fff00014fee01203fef01102;
assign testcases[409] = 512'hfef00012fef00012fff00123fff00122fff00012fff00012ede12213fed12313fef00003fef00003fff00003fff00003fff00005fff00014fee01203ede02202;
assign testcases[410] = 512'hfef00112fef00012ffe00223fff00123fef00112fef00112edd23313edd13314fef00004fef00003fff00003fff00003fff00005fff00014fed02304ede12203;
assign testcases[411] = 512'hfef00112fef00112ffe00223ffe00223fef00113fef00112edd23314edc23414fef00004fef00104fff00003fff00003fff00005fff00014fed02304ede13303;
assign testcases[412] = 512'hfef00122fef00122ffe00223ffe00233fef00123fef00112edd24414fdc24414fef00104fef00104ffe00004fff00003fff00005fff00015fed02404fde13303;
assign testcases[413] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef01113ecd24424edc24425fef00104fef00104ffe00004fff00003fff00005fff00025fec02405edd13304;
assign testcases[414] = 512'hfef00122fef01122ffe00233ffe01233fef01123fef01113edd24424edc25525fef00104fef00104ffe00104fff00003fff00005fff00025fec03405edd14404;
assign testcases[415] = 512'hfef00123fef01122ffe00233ffe01233fef01123fef01113edc35525fdc25525fef00104fef00104ffe00104fff00103fff00005fff00025fec13505fdd14404;
assign testcases[416] = 512'hfef00123fef01122ffe00234ffe01233fef01123fef01113edc35525edb25525fef00104fef00104ffe00104fff00103fff00005fff00025fec13505edd14404;
assign testcases[417] = 512'hfef00123fef01122ffe00234ffe01234fef01123fef01113edc35525edb25526fef00104fef00104ffe00104fff00103fff00005fff00025fdc13505edd14404;
assign testcases[418] = 512'hfef00123fef01122ffd01334ffd01234fef01123fef01113ecc35525ecb36626fef00104fef00104ffe00104fff00104fff00015fff00025edc13506ecd15404;
assign testcases[419] = 512'hfdf00123fef01122ffd01234ffd01234fef01133fef01123ecc35525ecb36626fef00104fef00104ffe00104fff00104fff00015fff00025fdb13506ecd15405;
assign testcases[420] = 512'hfef00123fef01122ffd01334ffd01234fef01123fef01123ecc36625fdb36626fef00104fef00104ffe00104fff00104fff00015fff00125feb14606edd15505;
assign testcases[421] = 512'hfef00123fef01122ffd01334ffd01344fef01123fef01123ecc36625fdb37626fef00104fef00104ffd00104fff00104fff00015fff00125feb14606fdd15505;
assign testcases[422] = 512'hfef00012fef00001fff00112fff00012fff00012fff00002fef11101fff11102fef00003fef00003fff00002fff00002fff00004fff00014fff01102fef11101;
assign testcases[423] = 512'hfef00012fef00012fff00122fff00122fff00012fff00012eee11212fee11213fef00003fef00003fff00003fff00002fff00005fff00014fee01203fef01102;
assign testcases[424] = 512'hfef00012fef00012fff00123fff00122fff00012fff00012ede12213fed12313fef00003fef00003fff00003fff00002fff00005fff00014fee01303ede02202;
assign testcases[425] = 512'hfef00112fef00012fff00223fff00123fef00112fff00012edd23313edd13314fef00003fef00003fff00003fff00003fff00005fff00014fed02304ede12203;
assign testcases[426] = 512'hfef00122fef00112ffe00223ffe00223fef00113fef00112edd23314edc24414fef00004fef00104fff00003fff00003fff00005fff00014fed02304fde13303;
assign testcases[427] = 512'hfef00122fef00122ffe00233ffe00233fef00123fef00112fdd23424fdc24425fef00104fef00104ffe00004fff00003fff00005fff00025fed02404fde13303;
assign testcases[428] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef00112ecd24414edc24415fef00104fef00104ffe00004fff00003fff00005fff00015eec02405edd13304;
assign testcases[429] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef01113edd24414edc25515fef00104fef00104ffe00004fff00003fff00005fff00025eec03405edd14404;
assign testcases[430] = 512'hfef00122fef01122ffe00233ffe00233fef01123fef01113edc24425edb25525fef00104fef00104ffe00004fff00003fff00005fff00025fdc03505edd14404;
assign testcases[431] = 512'hfef00122fef01122ffe00234ffe01233fef01123fef01113edc35525edb25526fef00104fef00104ffe00104fff00003fff00005fff00025eec03505edd14404;
assign testcases[432] = 512'hfef00133fef01132ffe01334ffe01234fef01133fef01123edc35525fdb26526fef00104fef00104ffe00104fff00103fff00015fff00025fec13506fdd14404;
assign testcases[433] = 512'hfef00123fef01122ffd01334ffe01234fef01123fef01123ecc35525edb36626fef00104fef00104ffe00104fff00103fff00015fff00025fdc13506ecd15404;
assign testcases[434] = 512'hfdf00123fef01122ffd01234ffd01234fef01123fef01123ecc35525edb25626fef00104fef00104ffe00104fff00104fff00015fff00025eec13506edd14405;
assign testcases[435] = 512'hfef00123fef01122ffd01334ffd01244fef01123fef01123ecc36625fdb36626fef00104fef00104ffd00104fff00104fff00015fff00125fdb14606ecd15505;
assign testcases[436] = 512'hfef00002fef00001fff00112fff00012fff00002fff00002fef11101fff01102fef00003fef00003fff00002fff00002fff00004fff00014fff01102fef01101;
assign testcases[437] = 512'hfef00012fef00012fff00122fff00122fff00012fff00012ede12213fed12313fef00003fef00003fff00003fff00002fff00005fff00014fed01203ede02203;
assign testcases[438] = 512'hfef00112fef00012fff00223fff00123fff00112fff00012edd23313fed13314fef00003fef00003fff00003fff00003fff00005fff00014fed02304ede12203;
assign testcases[439] = 512'hfef00012fef00011fff00112fff00012fff00012fff00002fef01112fff01112fef00003fef00003fff00003fff00002fff00004fff00014fff00102fef01102;
assign testcases[440] = 512'hfef00012fef00012fff00122fff00122fff00012fff00012fee12212fee12213fef00003fef00003fff00003fff00002fff00005fff00014fee01203fef01102;
assign testcases[441] = 512'hfef00012fef00012fff00123fff00122fff00012fff00012ede12313fed12313fef00003fef00003fff00003fff00003fff00005fff00014fed01303fde02203;
assign testcases[442] = 512'hfef00112fef00012ffe00223fff00123fef00112fff00112edd23313fdd13314fef00003fef00003fff00003fff00003fff00005fff00014fed02304ede12203;
assign testcases[443] = 512'hfef00122fef00112ffe00223ffe00223fef00123fef00112edd23314edc24414fef00004fef00104fff00003fff00003fff00005fff00014fed02304fde13303;
assign testcases[444] = 512'hfef00122fef00122ffe00233ffe00233fef01123fef01112edd25424fdc25425fef00104fef00104ffe00004fff00003fff00005fff00015fec03405edd14304;
assign testcases[445] = 512'hfef00112fef00012fff00123fff00123fff00112fef00112fff00101fff00001fef00003fef00003fff00003fff00003fff00005fff00014fff00001fef00001;
assign testcases[446] = 512'hfef00112fef01112ffe01333ffe01233fef01113fef01113fef11112fff01111fef00104fef00104ffe00104fff00103fff00005fff00015fff01102fef01101;
assign testcases[447] = 512'hfef10122fef01122ffd01334ffd01334fef01123fef01113ede12212fee11212fef00104fef00104ffd00105fff00104fff00005fff00125fee01202fee01102;
assign testcases[448] = 512'hfef10223fef01123ffd01444ffd01344fef01123fef11223fde12312fee12212fef01104fef01104ffd00105fff00104fff00015fff00125fee01202fde02202;
assign testcases[449] = 512'hfdf10223fef01223ffc01445ffd01445fef01223fef11223fdd12213fee12212fef01104fef01104ffd00106fff00105fff00016fff00125fee01203fde02202;
assign testcases[450] = 512'hfde11233fde12233ffb02556ffc01456fee12234fee12224fdd23323fed13313fde11205fde01205ffc01106fff01105fff00016ffe00136fed02303fde12203;
assign testcases[451] = 512'hfde11334fde12234fea02656ffb02566fde12234fee12234ecc24424fdc23423fde11205fde11205ffb01107fff01106fff00016ffe00136fed02303fdd13303;
assign testcases[452] = 512'hfce11344fde12344fea02667ffa02567fdd13344fde12334ecc35424fdc24424fdd11206fdd11206ffa01108ffe01107fff00017fed00136fec02404fcd13303;
assign testcases[453] = 512'hfcd21345fcd13344fe902778fea02677fdd13345fdd13335ecb35525fdb24424fdd11206fdd11306fea01208ffe01107fff00017fed00147fec03404fcc14404;
assign testcases[454] = 512'hfcd21455fcd13455fe802778fe902688fdd13345fdd13445ebb36535fcb25525fcd11306fcc11307fe901209ffe01208ffe00017fec00247fdc03504ecc14404;
assign testcases[455] = 512'hfcc21455fcc13455fe802779fe802789fcc13455fcc13445eba36635fcb25525fcc11307fcc11307fe80120affe01208ffe00018fec00247fdb13505ecc15404;
assign testcases[456] = 512'hfbc21556fbc13455fe702889fe813799fcc13456fcc13446eba46636fca36625fcc11307fcc11407fe80120affe01209ffe00118feb00258fdb13505ecc15505;
assign testcases[457] = 512'hfbc21566fbc14566fe70388afe71389afcc13456fcc14546ebad9736fca37625fbb11407fbb12408fe70120bffe01209ffe00118feb00258fdb14605ecb16505;
assign testcases[458] = 512'hfbb21566fbb14566fe60289afe7138aafcb13566fcb14556eb947736fca37636fbb11408fbb12408fe60120bffd0120affe00118feb00258fdb14605ebb16605;
assign testcases[459] = 512'hfef00112fef01112fff00223fff00223fff00112fff00112fff00101fff00001fef00103fef00103fff00003fff00003fff00005fff00014fff00001fef00001;
assign testcases[460] = 512'hfef00112fef01112ffe01333ffe01233fef01113fef01113fef11112fff01111fef00104fef00104ffe00104fff00103fff00005fff00015fff00102fef01101;
assign testcases[461] = 512'hfef10123fef01122ffd01334ffd01334fef01123fef01113fee11212fee11112fef00104fef00104ffe00105fff00104fff00005fff00125fff01102fef01102;
assign testcases[462] = 512'hfdf10223fdf01223ffd01445ffd01344fef01123fef11223ede12212fee12212fef01104fef01104ffd00105fff00104fff00016fff00125fee01202fde01102;
assign testcases[463] = 512'hfdf10223fdf02223ffc01445ffd01445fef01223fef12223fdd12323fee12212fef01105fef01205ffd00106fff00105fff00016ffe00125fee01203fde02202;
assign testcases[464] = 512'hfde11234fde12233ffb01556ffc01556fee12234fde12224edd23323fed13323fde11205fde01205ffc01107fff01106fff00016ffe00136fed02303ede12203;
assign testcases[465] = 512'hfde11334fde12334ffa02657ffb02566fde12334fde12334ecc24424fdc23424fde11205fde11206ffb01107fff01106fff00016ffd00136fed02304fdd13303;
assign testcases[466] = 512'hfcd11344fdd13344fea02667fea02667fdd12345fdd13335ecb34424fdc24424fdd11206fdd11306ffa01108ffe01107fff00017fed00137fec02404fcd13303;
assign testcases[467] = 512'hfcd21445fcd13345fe902778fe902678fdd13345fdd13335ecb35535fdb25424fcd11306fdd11306fe901209ffe01207fff00017fed00247fec03404fcc14404;
assign testcases[468] = 512'hfcd21455fcd13455fe802778fe902788fdd13445fdd13445ebb36535fdb25525fcc11307fcc11307fe901209ffe01208ffe00017fec00247fdc03504fcc14404;
assign testcases[469] = 512'hfcc21555fcc13455fe802779fe812789fdc13456fcc13446eba36635fcb25525fcc11307fcc11407fe80120affe01208ffe00118fec00248fdb13505ecc15404;
assign testcases[470] = 512'hfbc21556fbc14556fe702889fe813799fcc13456fcc14446eba46636fca36635fcc11407fcc12407fe70120affe01209ffe00118feb00258fdb13505ecc15505;
assign testcases[471] = 512'hfbb21566fbb14566fe60388afe71389afcb13566fcb24556eba47736fca36636fbb11408fbb12408fe70120bffe01209ffe00118feb01258fdb14605ecb15505;
assign testcases[472] = 512'hfbb21666fbb14566fe60389afe7138aafcb13566fcb24557eb947736fca37636fbb11408fbb12408fe60120bffd0120affe00129fea01258fdb14605ebb16505;
assign testcases[473] = 512'hfef00112fef00112fff00123fff00123fff00112fff00112fff00101fff00001fef00004fef00003fff00003fff00003fff00005fff00014fff00001fef00001;
assign testcases[474] = 512'hfef00122fef01112ffe01234ffe01233fef01113fef01113fef11112fff01111fef00104fef00104ffe00104fff00103fff00005fff00015fff00102fef01101;
assign testcases[475] = 512'hfef10123fef01122ffd01334ffd01334fef01123fef01113fee11212fee11112fef00104fef00104ffd00105fff00104fff00005fff00125fff01102fef01102;
assign testcases[476] = 512'hfef10223fef01223ffd01445ffd01344fef01223fef11223fde12222fee12212fef01104fef01104ffd00105fff00104fff00016fff00125fee01202fee01102;
assign testcases[477] = 512'hfdf10223fdf02223ffc01445ffd01445fee02223fef12223fdd12323fee12212fef01105fee01205ffd00106fff00105fff00016ffe00125fee01203fde02202;
assign testcases[478] = 512'hfde11334fde12233ffb01556ffc01556fee12234fee12224fdd23323fed13323fde11205fde01205ffc01107fff01106fff00016ffe00136fed02303fde12203;
assign testcases[479] = 512'hfde11344fde12344ffa02667feb02566fde12334fde12334ecc24434fdc23424fde11206fdd11206ffb01107fff01106fff00017fed00136fed02304fdd13303;
assign testcases[480] = 512'hfcd11344fcd13344fea02667fea02677fdd13345fdd13335ecc35534fdc24424fdd11206fdd11306ffa01208ffe01107fff00017fed00147fec02404fcd13304;
assign testcases[481] = 512'hfcd21445fcd13455fe902778fe902678fdd13345fdd13435ecb35535fdb25524fcd11306fcd11306fe901209ffe01207fff00017fec00247fec03404fcc14404;
assign testcases[482] = 512'hfcd21455fcd13455fe802778fe902788fdc13455fdd13445ebb36635fdb25535fcc11307fcc11307fe901209ffe01208ffe00118fec00247fdb03505fcc14404;
assign testcases[483] = 512'hfbc21556fcc14455fe802889fe813789fcc13456fcc14446eba36646fcb25535fcc11307fcc11407fe80120affe01209ffe00118fec00258fdb13505ecc15504;
assign testcases[484] = 512'hfbc21556fbc14566fe702889fe813799fcc13456fcc14546eba47646fca36635fcc11407fcb12407fe70120affe01209ffe00118feb01258fdb13505ecb15505;
assign testcases[485] = 512'hfbb21566fbb14566fe60288afe71389afcb14566fcb24556eba47746fca36636fbb12408fbb12408fe70120bffe01209ffe00118feb01258fdb14605ecb15505;
assign testcases[486] = 512'hfbb21667fbb14566fe60399afe6138aafcb14567fcb24557ea947746fca37636fbb12408fbb12508fe60120bffd0120affe00129fea01269fda14606ebb16505;
assign testcases[487] = 512'hfef00112fef00112fff00212fff00112fff00112fff00102fff00111fff00011fef00003fef00103fff00003fff00002fff00005fff00014fff00001fef00001;
assign testcases[488] = 512'hfef00122fef01122ffe01234ffe01233fef01113fef01113fef11112fff01111fef00104fef00104ffe00104fff00103fff00005fff00015fff00102fef01101;
assign testcases[489] = 512'hfef10123fef01123ffd01334ffd01334fef01123fef01113fee12212fee11112fef00104fef00104ffd00105fff00104fff00005fff00125fff01102fef01102;
assign testcases[490] = 512'hfdf10223fef01223ffd01445ffd01344fef01223fef11223fde12222fee12212fef01104fef01104ffd00105fff00104fff00016fff00125fee01202fee01102;
assign testcases[491] = 512'hfdf10223fdf02233ffc01445ffd01455fef02223fef12223fdd12323fee12222fef01105fde01205ffd00106fff00105fff00016ffe00125fee01203fde02202;
assign testcases[492] = 512'hfde11334fde12233ffb01556ffc01556fee12234fee12224fdd23323fed13323fde11205fde01205ffc01107fff01106fff00016ffe00136fed02303fde12203;
assign testcases[493] = 512'hfde11334fde12344ffa02657ffb02566fde12334fde12334ecc24434fdc23424fde11206fdd11206ffb01107fff01106fff00017fed00136fed02304fdd13303;
assign testcases[494] = 512'hfcd11344fcd13344fe902667fea02677fdd13345fdd13335ecc35534fdc24424fdd11206fdd11306ffa01108ffe01107fff00017fed00147fec02404fcd13304;
assign testcases[495] = 512'hfcd21445fcd13455fe902778fe902678fdd13345fdd13435ecb35535fdb25534fcd11306fcd11306fe901209ffe01207fff00017fec00247fec03404fcc14404;
assign testcases[496] = 512'hfcc21455fcd13455fe802778fe902788fdc13455fdc13445ebb36635fdb25535fcc11307fcc11307fe901209ffe01208ffe00118fec00247fdc03505fcc14404;
assign testcases[497] = 512'hfcc21556fcc14455fe802889fe813789fcc13456fcc14446eba46646fcb26535fcc11307fcc12407fe80120affe01209ffe00118fec00258fdb13505ecc15504;
assign testcases[498] = 512'hfbc21556fbc14566fe702889fe713899fcc13456fcc24546eba47646fca36635fcb12407fcb12408fe70120affe01209ffe00118feb01258fdb13505ecc15505;
assign testcases[499] = 512'hfbb21566fbb14566fe60288afe71389afcb14566fcb24556eba47746fca36636fbb12408fbb12408fe70120bffe01209ffe00118feb01258fdb14605ebb15505;
assign testcases[500] = 512'hfbb21667fbb14576fe60299afe6138aafcb14567fcb24557ea947746fca37636fbb12408fbb12508fe60120bffd0120affe00129fea01269fda14606ebb16505;
assign testcases[501] = 512'hfef00112fef00112fff00223fff00123fff00112fff00112fff00111fff00001fef00004fef00104fff00003fff00003fff00005fff00014fff00001fef00001;
assign testcases[502] = 512'hfef00122fef01122ffe01334ffe01233fef01113fef01113fef11112fff01111fef00104fef00104ffe00104fff00104fff00005fff00015fff00102fef01101;
assign testcases[503] = 512'hfef10223fef01123ffd01334ffd01334fef01123fef01113fee11212fee11112fef00104fef00104ffd00105fff00104fff00005fff00125fff01102fef01102;
assign testcases[504] = 512'hfdf10223fdf01223ffd01445ffd01344fef01223fef11223fde12222fee12212fef01104fef01104ffd00105fff00104fff00016fff00125ffe01202fee01102;
assign testcases[505] = 512'hfde10233fdf12233ffc01445ffc01445fee02224fef12223fdd12323fee12222fde01105fde01205ffc00106fff00105fff00016ffe00126fee01203fde02202;
assign testcases[506] = 512'hfde11334fde12234ffb01556ffb02556fde12234fde12224fcd23333fdd13323fde11205fde01205ffb01107fff01106fff00016fee00136fed02303fde12203;
assign testcases[507] = 512'hfde11344fde13344ffa02667feb02567fde12334fde12334ecc24434fdc23424fdd11206fdd11206ffb01107fff01106fff00017fed00136fed02304fdd13303;
assign testcases[508] = 512'hfcd11445fcd13344fe902667fea02677fdd13345fdd13335ecc35534fdc24434fdd11306fdd11306ffa01208ffe01107fff00017fed00247fec02404fdd13304;
assign testcases[509] = 512'hfcd21445fcd13455fe902778fe902678fdd13345fdd13435ecb35535fdb25534fcd11306fcc11307fe901209ffe01208ffe00017fec00247fdc03404ecc14404;
assign testcases[510] = 512'hfcc21455fcc13455fe802779fe902788fdc13455fdc13445ebb36645fdb25535fcc11307fcc11407fe901209ffe01208ffe00118fec00247fdc03505ecc14404;
assign testcases[511] = 512'hfcc21556fcc14556fe802889fe813789fcc13456fcc14446eba36646fcb25535fcc11307fcc12407fe80120affe01209ffe00118feb00258fdb13505ecc15504;
assign testcases[512] = 512'hfbc21556fbc14566fe603889fe71389afcb14456fcc24546eba47646fca36635fcb12408fbb12408fe70120bffe01209ffe00118feb01258fdb13505ecc15505;
assign testcases[513] = 512'hfbb21666fbb14566fe61398afe71389afcb14566fcb24546eba47736fca36636fbb12408fbb12408fe70120bffd0120affe00119feb01258fdb13605ebb16505;
assign testcases[514] = 512'hfab21667fbb14667fe51399afe71389bfcb14567fcb24557da948736eca37636fbb12408fbb12508fe60120cffd0120affe00119fea01259eda14605ebb16605;
assign testcases[515] = 512'hfcd21455fcd14464ffb01455ffc01455fcc14565fcc24556fff00000fff00001fcc12406fcc12406ffb01106fff01105ffe00128feb01368fff00001fef00001;
assign testcases[516] = 512'hfcd21565fcd14565ffa01566ffb01465fcb14576fcc25656fff00000fff00001fcc12407fcc12407ffb01107fff01106ffe00129fea01368fff00001fef00001;
assign testcases[517] = 512'hfcc21565fcc25575fea01566feb02566fcb15676fcb25666fff00001fff00001fcc12407fcc12507fea01107ffe01106ffd00129fda01379fff00001fef00001;
assign testcases[518] = 512'hfbc21676fbc25675fea02667fea02576fba15687fbb26767fff00001fff00001fbb22508fbb12508fea01108ffe01107ffd00129fd901489fff00101fef00001;
assign testcases[519] = 512'hfbc32676fbc26686fe902677fea02577fba26787fba36777fff00001fff00001fbb22508fbb13608fe901208ffe01107ffd0012afd80148afff00101fef00001;
assign testcases[520] = 512'hfbb32786fbb26686fe802677fe902687fb926798fba37878fff00001fff00001fba23508fba13608fe901208ffe01207ffd0112afd80148afff00101fef00001;
assign testcases[521] = 512'hfef00112fef00112fff00112fff00112fef00113fef00112fff00000fff00000fef00104fef00104fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[522] = 512'hfef00122fef01122ffe00223fff00123fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00015fff00125fff00001fff00000;
assign testcases[523] = 512'hfef10223fdf01233ffe00233ffe00233fef01233fef11223fff00000fff00000fef01104fef01204ffe00104fff00103fff00016ffe00136fff00001fff00001;
assign testcases[524] = 512'hfdf10233fdf12233ffe01234ffe01233fee02234fee12234fff00000fff00000fde01205fde01205ffe00104fff00104fff00016ffe00136fff00001fef00001;
assign testcases[525] = 512'hfde11333fde12233ffd01334ffe01234fee12344fde12334fff00000fff00000fde11205fde01205ffd00105fff00104fff00016fed00236fff00001fef00001;
assign testcases[526] = 512'hfde11344fde13344ffc01344ffd01344fdd13445fdd13445fff00000fff00000fdd11306fdd11306ffd00105fff00105fff00117fec00247fff00001fef00001;
assign testcases[527] = 512'hfcd31454fcd24454ffc01455ffc01455fdd24455fdd34545fff00000fff00000fcd22306fdd22406ffc00106fff00105ffe00118fec01257fff00001fef00001;
assign testcases[528] = 512'hfcd21555fcd14454ffb01555ffc01455fcc14566fcc24556fff00000fff00001fcc12407fcc12407ffb01106fff00105ffe00128feb01368fff00001fef00001;
assign testcases[529] = 512'hfcd21565fcd15565ffb01566ffb01466fcb14566fcb25656fff00000fff00001fcc12407fcc12407ffb01107fff01106ffe00129fea01369fff00001fef00001;
assign testcases[530] = 512'hfcc21565fcc25575fea01566feb02576fcb15677fcb26767fff00001fff00001fcb12507fcc12507fea01107ffe01106ffd00129fda01379fff00001fef00001;
assign testcases[531] = 512'hfbc31676fbc26676fe902677fea02576fba15787fba26767fff00001fff00001fbb22508fbb12508fe901108ffe01107ffd0012afd90147afff00001fef00001;
assign testcases[532] = 512'hfbc32676fbc26676fe902677fea02577fba26787fba37877fff00001fff00001fbb23508fbb13608fe901208ffe01207ffd0012afd80148afff00101fef00001;
assign testcases[533] = 512'hfbb32776fbb26786fe802678fe902687fb926798fb937878fff00011fff00011fba23608fba13608fe901209ffe01207ffd0112afd80148afff00101fef00001;
assign testcases[534] = 512'hfef00112fef00112fff00112fff00112fef00113fef00112fff00000fff00000fef00104fef00104fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[535] = 512'hfef00122fef01122ffe00223fff00123fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00015fff00125fff00001fff00000;
assign testcases[536] = 512'hfef10223fdf01223ffe00233ffe00233fef01223fef11223fff00000fff00000fef01104fef01204ffe00104fff00103fff00016ffe00126fff00001fff00001;
assign testcases[537] = 512'hfdf10233fdf12233ffe01333ffe01233fee02234fee12224fff00000fff00000fde01205fde01205ffe00104fff00104fff00016ffe00136fff00001fef00001;
assign testcases[538] = 512'hfde11333fde12233ffd01334ffe01234fee12334fde12334fff00000fff00000fde11205fde01205ffd00105fff00104fff00016fed00136fff00001fef00001;
assign testcases[539] = 512'hfde11344fde13344ffc01444ffd01344fdd13445fdd13435fff00000fff00000fdd11306fdd11306ffd00105fff00104fff00117fed00247fff00001fef00001;
assign testcases[540] = 512'hfcd21444fcd13454ffc01445ffc01455fdd13455fdd14545fff00000fff00000fcd11306fdd12406ffc00106fff00105ffe00118fec01257fff00001fef00001;
assign testcases[541] = 512'hfcd21555fcd14454ffb01555ffc01455fcc14566fcc24556fff00000fff00001fcc12406fcc12407ffb01106fff00105ffe00128feb01358fff00001fef00001;
assign testcases[542] = 512'hfcd21555fcd25565ffa01556ffb01466fcb14566fcb25656fff00000fff00001fcc12407fcc12507ffb01107fff01106ffe00129fea01369fff00001fef00001;
assign testcases[543] = 512'hfcc21565fcc25565fea01566feb02566fcb15677fcb26767fff00000fff00001fcb12507fcb12507fea01107ffe01106ffd00129fda01379fff00001fef00001;
assign testcases[544] = 512'hfbc21666fbc26675fe902667fea02576fba15677fba26767fff00001fff00001fbb22508fbb12508fea01108ffe01107ffd0012afd901479fff00001fef00001;
assign testcases[545] = 512'hfbc32676fbc26676fe902677fea02577fba26787fba37867fff00011fff00001fbb23508fbb13608fe901208ffe01207ffd0012afd80148afff00101fef00001;
assign testcases[546] = 512'hfbb32776fbb26786fe802678fe902687fb926788fb937878fff00011fff00011fba23608fba13608fe801209ffe01208ffc0112afd80148afff00101fef00001;
assign testcases[547] = 512'hfbb32787fbb27786fe802788fe902688fa926898fa937978fff00011fff00111fba23609fba13609fe801209ffe01208ffc0112bfd70149bfff00101fef00001;
assign testcases[548] = 512'hfab32776fbb26786fe802788fe902688fa926888fb937878fff00001fff00011fba23609fba13608fe801209ffe01208ffc0112bfd80148afff00101fef00001;
assign testcases[549] = 512'hfab32756fbb27766fe802767fe902667fb927868fb937858fff00011fff00011fba23608fba23608fe801209ffe01207ffc0112afd80146afff00101fef00001;
assign testcases[550] = 512'hfab21866fbb25867fe713968fe913878fa915888fa925968fff46601fff36501fba12609fba12708fe801209ffe01208ffc0012bfd70148bfff13501fef15401;
assign testcases[551] = 512'heab42766ebb27767fe802778fe902678fa927888fa938968fff00101fff00101eba23609eba23608fe801209ffe01208ffc0112bfd70157bfff00101fef00001;
assign testcases[552] = 512'hfde11333fde12333ffd01334ffe01334fee12334fde12334fff00000fff00000fde11205fde01205ffd00105fff00104fff00017fed00236fff00001fef00001;
assign testcases[553] = 512'hfde11333fde12333ffd01334ffe01234fee12334fde12334fff00000fff00000fde11205fde01205ffd00105fff00104fff00017fed00236fff00001fef00001;
assign testcases[554] = 512'hfde21323fde22323ffd01324ffe11323fde12324fde12324fff00000fff00000fde11205fde11305ffd00104fff00104fff00017fed00226fff00001fef00001;
assign testcases[555] = 512'hfde11333fde12333ffd01334ffd01234fde12334fde12324fff00000fff00000fde11205fde11205ffd00105fff00104fff00017fed00236fff00001fef00001;
assign testcases[556] = 512'hfde11333fde12333ffd01334ffe01234fde12334fde12334fff00000fff00000fde11205fde11305ffd00105fff00104fff00017fed00236fff00001fef00001;
assign testcases[557] = 512'hfde11333fde12333ffd01334ffd01334fde12334fde13334fff00000fff00000fde11205fde11305ffd00105fff00104fff00017fed00236fff00001fef00001;
assign testcases[558] = 512'hfab32777fab38787fe802788fe902688ea927898da938978fff00011fff00111eaa23609faa23609fe801209ffe01208ffc0112bfc70158bfff00101fef00001;
assign testcases[559] = 512'hfbb32777fbb37777fe802788fe802688fa927888fa938978fff00011fff00001fba23609fba23609fe801209ffe01208ffc0112bfd70158bfff00101fef00001;
assign testcases[560] = 512'hfbb32787fbb27787fe802788fe902688fa927898fa938988fff00011fff00011fba23609fba23609fe801209ffe01208ffc0113bfd70159bfff00101fef00001;
assign testcases[561] = 512'hfbb32777fbb27787fe802788fe802688fa927889fa938978fff00001fff00001fba23609fba23609fe801209ffe01208ffc0112bfd70158bfff00001fef00001;
assign testcases[562] = 512'hfbc32676fbb27676fe902677fe902677fba26788fba37868fff00000fff00001fbb23508fbb13608fe901209ffe01208ffd0112afd80148afff00001fef00001;
assign testcases[563] = 512'hfbc32666fbb27676fe902677fe902577fba26788fba37868fff00000fff00001fbb23508fbb13608fe901209ffe01207ffd0112afd80147afff00001fef00001;
assign testcases[564] = 512'hfab217b6fbb157c7fe802888fe902798fb9147c8fb9258a8fef59811fff4a912fba12508fba12608fe801209ffe01208ffd0013afd8014bafff16902fef29701;
assign testcases[565] = 512'hfab32786fbb26796fe802778fe902688fb9167a8fb937888fff12211fff12211fba22508fba13608fe801209ffe01208ffd0013afd80149afff01201fef01201;
assign testcases[566] = 512'hfef00112fef01112fff00112fff00112fff01112fef01112fff00000fff00000fef00104fef00104fff00003fff00002fff00005fff00015fff00001fff00001;
assign testcases[567] = 512'hfef10122fef01122fff01223fff01222fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00015fff00125fff00001fff00001;
assign testcases[568] = 512'hfef10233fef01233ffe01223ffe01233fef01233fef11223fff00001fff00001fef01104fef01104ffe00104fff00103fff00016fff00135fff00001fef00001;
assign testcases[569] = 512'hfdf10233fdf02233ffe01233ffe01233fee02233fee12234fff00001fff00001fdf01205fef01204ffe00104fff00103fff00016ffe00136fff00001fef00001;
assign testcases[570] = 512'hfde11233fde12233ffd01334ffe01234fee12234fee12334fff00001fff00001fde11205fde01205ffe00105fff00104fff00016ffe00136fff00001fef00001;
assign testcases[571] = 512'hfde11344fde13344ffd01344ffd01344fdd13344fdd13435fff00001fff00101fde11305fde11305ffd00105fff00104fff00017fed00247fff00101fef00001;
assign testcases[572] = 512'hfcd21454fcd13454ffc01445ffc01355fdd13455fdd14545fff00001fff00101fdd11306fdd11306ffc00106fff00105ffe00117fec01257fff00101fef00001;
assign testcases[573] = 512'hfcd21455fcd14455ffb01455ffc01455fcc14565fcc24546fff00001fff00001fcd12406fcd12406ffb01106fff01105ffe00118feb01258fff00001fef00001;
assign testcases[574] = 512'hfcd21565fcd14565ffb01556ffb01456fcc14566fcc25656fff00001fff00001fcc12407fcc12407ffb01107fff01106ffe00128feb01368fff00001fef00001;
assign testcases[575] = 512'hfcc21565fcc25565fea01556ffb01466fcb14576fcb25656fff00001fff00001fcc12407fcc12407ffb01107fff01106ffe00129fea01368fff00001fef00001;
assign testcases[576] = 512'hfbc21575fcc25575fea02566feb01566fcb15686fcb25666fff00001fff00101fcc12407fcc12507ffa01107ffe01106ffd00129fda01379fff00001fef00001;
assign testcases[577] = 512'hfbc21676fbc25686fe902577fea02577fba15687fbb26777fff00001fff00101fbb12508fbb12507fea01108ffe01107ffd00129fd901389fff00101fef00001;
assign testcases[578] = 512'hfbc32686fbc26686fe902677fea02577fba15797fba26777fff00001fff00101fbb22508fbb12508fe901208ffe01107ffd0012afd901489fff00101fef00001;
assign testcases[579] = 512'hfbb32686fbb26696fe802677fe902687fba15797fba26878fff12211fff12211fba22508fbb12508fe901208ffe01207ffd0012afd80149afff01201fef02201;
assign testcases[580] = 512'hfef00112fef01112fff00112fff00112fef01112fef01112fff00000fff00000fef00104fef00104fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[581] = 512'hfef00122fef01122fff00223fff00123fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00015fff00125fff00001fff00000;
assign testcases[582] = 512'hfef10233fef01233ffe01223ffe01233fef01233fef11223fff00000fff00000fef01104fef01104ffe00104fff00103fff00016ffe00135fff00001fff00001;
assign testcases[583] = 512'hfdf10233fdf12233ffe01233ffe01233fee02234fee12234fff00000fff00000fde01205fde01205ffe00104fff00103fff00016ffe00136fff00001fef00001;
assign testcases[584] = 512'hfde11233fde12233ffd01334ffe01234fee12344fee12334fff00000fff00001fde11205fde01205ffe00105fff00104fff00016ffe00146fff00001fef00001;
assign testcases[585] = 512'hfde11344fde13344ffd01344ffd01344fdd13344fdd13434fff00001fff00001fde11305fde11305ffd00105fff00104fff00117fed00246fff00001fef00001;
assign testcases[586] = 512'hfde11454fde13454ffc01445ffd01355fdd13455fdd13445fff00001fff00001fdd11306fdd11306ffc00106fff00105ffe00117fec00257fff00001fef00001;
assign testcases[587] = 512'hfcd21454fcd14464ffc01455ffc01455fdc14465fcc24555fff00001fff00001fcd11306fcd12406ffc00106fff00105ffe00128fec01267fff00001fef00001;
assign testcases[588] = 512'hfcd21465fcd14465ffb01456ffc01465fcc14576fcc24556fff00001fff00001fcc12407fcc12406ffb01106fff01106ffe00128feb01368fff00001fef00001;
assign testcases[589] = 512'hfcd21565fcd15575fea01566ffb01466fcb14576fcb25666fff00001fff00001fcc12407fcc12407ffb01107fff01106ffe00129feb01378fff00001fef00001;
assign testcases[590] = 512'hfbc21575fcc25575fea02566feb01576fcb15686fcb25667fff00001fff00001fcc12407fcc12507ffa01107ffe01106ffd00129fda01389fff00001fef00001;
assign testcases[591] = 512'hfbc21686fbc25686fe902577fea02577fba15697fba26777fff00001fff00001fbb12508fbb12507fea01108ffe01107ffd00129fd901389fff00001fef00001;
assign testcases[592] = 512'hfbb32686fbb26686fe902677fea02577fba16797fba26777fff00001fff00001fbb22508fbb12508fe901208ffe01107ffd0012afd901499fff00001fef00001;
assign testcases[593] = 512'hfbb32786fbb26696fe802778fe902687fb9267a8fb936888fff12211fff12211fba22508fba13608fe901209ffe01208ffd0013afd80149afff01201fef02201;
assign testcases[594] = 512'hfef00112fef01112fff00112fff00112fef01113fef01112fff00000fff00000fef00104fef00104fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[595] = 512'hfef00122fef01122fff00223fff00123fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00015fff00125fff00001fff00000;
assign testcases[596] = 512'hfef10233fef01233ffe01223ffe01233fef01233fef11223fff00000fff00000fef01104fef01104ffe00104fff00103fff00016ffe00135fff00001fff00001;
assign testcases[597] = 512'hfdf10233fdf12233ffe01233ffe01233fee02234fee12234fff00000fff00000fde01205fde01205ffe00104fff00103fff00016ffe00136fff00001fff00001;
assign testcases[598] = 512'hfde11233fde12233ffd01334ffe01233fee12334fee12334fff00000fff00000fde11205fde01205ffe00104fff00104fff00016ffe00136fff00001fef00001;
assign testcases[599] = 512'hfde11344fde13344ffd01344ffd01344fdd13344fdd13434fff00000fff00001fde11205fde11305ffd00105fff00104fff00017fed00246fff00001fef00001;
assign testcases[600] = 512'hfde11444fde13454ffc01445ffd01345fdd13455fdd13445fff00000fff00001fdd11306fdd11306ffc00106fff00105ffe00117fec01257fff00001fef00001;
assign testcases[601] = 512'hfcd21454fcd14454ffc01455ffc01455fdc14465fcc24545fff00000fff00001fcd12306fcd12406ffc00106fff00105ffe00118fec01257fff00001fef00001;
assign testcases[602] = 512'hfcd21565fcd14465ffb01456ffc01455fcc14566fcc24556fff00001fff00001fcc12407fcc12406ffb01107fff01106ffe00128feb01368fff00001fef00001;
assign testcases[603] = 512'hfcd21565fcd15565fea01566ffb01466fcb14576fcb25656fff00001fff00001fcc12407fcc12407ffb01107fff01106ffe00128feb01368fff00001fef00001;
assign testcases[604] = 512'hfbc21565fbc25575fea02566feb01566fcb15676fcb25666fff00001fff00001fcc12407fcc12507ffa01107ffe01106ffd00129fda01379fff00001fef00001;
assign testcases[605] = 512'hfbc21676fbc25676fe902567fea02577fba15687fbb26767fff00001fff00001fbb12508fbb12507fea01108ffe01107ffd00129fd901379fff00001fef00001;
assign testcases[606] = 512'hfbc32686fbc26686fe902677fea02577fba15797fba26777fff00001fff00001fbb22508fbb12508fe901208ffe01107ffd0012afd901489fff00001fef00001;
assign testcases[607] = 512'hfbb32686fbb26686fe802677fe902687fb926798fba26878fff12211fff12211fba22508fbb12608fe901209ffe01207ffd0012afd80149afff01201fef01201;
assign testcases[608] = 512'hfbb327c6fbb266c6fe902787fea02797fba157d7fba267a7fff24411fff25511fbb12508fbb12508fe901208ffe01207ffd00139fd9014c9fff03501fef14401;
assign testcases[609] = 512'hfbb216a6fbb256a6fe901687fea01597fba156b7fba25797fff11101fff11111fbb12508fbb12508fe901108ffe01107ffd00139fd9013a9fff01101fef01101;
assign testcases[610] = 512'hfef00112fef01112fff00112fff00112fff01112fff00112fff00000fff00000fef00103fef00103fff00003fff00002fff00005fff00014fff00001fff00000;
assign testcases[611] = 512'hfef00122fef01122fff00122fff00122fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00002fff00015fff00025fff00001fff00000;
assign testcases[612] = 512'hfef10132fef01132ffe00233fff00133fef01133fef01123fff00000fff00000fef00104fef00104fff00004fff00003fff00015fff00135fff00001fff00001;
assign testcases[613] = 512'hfef10233fef01233ffe01233ffe01233fef01233fef11233fff00000fff00000fef01104fef01104ffe00104fff00103fff00016ffe00135fff00001fef00001;
assign testcases[614] = 512'hfdf10233fdf01243ffe01233ffe01233fee02243fee12233fff00000fff00000fdf01205fdf01204ffe00104fff00103fff00016ffe00135fff00001fef00001;
assign testcases[615] = 512'hfde11343fde12243ffd01344ffe01244fde12354fde12344fff00000fff00001fde11205fde01205ffd00105fff00104fff00016ffe00146fff00001fef00001;
assign testcases[616] = 512'hfde11354fde13354ffd01344ffd01354fdd13354fdd13444fff00001fff00001fde11205fde11305ffd00105fff00104fff00017fed00256fff00001fef00001;
assign testcases[617] = 512'hfce11464fde13364ffc01455ffd01355fdd13465fdd13455fff00001fff00001fdd11306fdd11306ffc00106fff00105ffe00127fec00267fff00001fef00001;
assign testcases[618] = 512'hfcd21474fcd13474ffb01465ffc01465fcc13475fcc14565fff00001fff00001fcd11306fcd11306ffc00106fff00105ffe00128fec01277fff00001fef00001;
assign testcases[619] = 512'hfcd21575fcd14475ffb01566ffb01466fcc14586fcc24566fff00001fff00001fcc12407fcc12407ffb01107fff01106ffe00128feb01388fff00001fef00001;
assign testcases[620] = 512'hfbc21575fcc25575fea01566feb01576fcb15686fcb25666fff00001fff00001fcc12407fcc12507ffa01107ffe01106ffd00129fda01388fff00001fef00001;
assign testcases[621] = 512'hfbc21686fbc25686fe902677fea02577fba15697fba26777fff00001fff00001fbb12508fbb12507fea01108ffe01107ffd00129fd901389fff00001fef00001;
assign testcases[622] = 512'hfbb32686fbb26696fe902677fea02587fba26797fba26777fff00001fff00001fbb22508fbb13508fe901208ffe01207ffd0012afd90149afff00001fef00001;
assign testcases[623] = 512'hfbb32796fbb26696fe802688fe902688fb9267a8fb926888fff11201fff12211fba22508fba12608fe901209ffe01208ffd0013afd8014aafff01201fef01101;
assign testcases[624] = 512'hfef00112fef01112fff00112fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[625] = 512'hfef00122fef01122fff00223fff00223fef01123fef01223fff00000fff00000fef00104fef00104fff00004fff00003fff00015fff00125fff00001fff00000;
assign testcases[626] = 512'hfef10233fef01233ffe01223ffe01233fef01233fef11223fff00000fff00000fef01105fef01204ffe00104fff00103fff00016ffe00135fff00001fff00001;
assign testcases[627] = 512'hfdf10233fdf12233ffe01333ffe01233fee02234fee12334fff00000fff00000fde01205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00001;
assign testcases[628] = 512'hfde11333fde12233ffd01334ffe01234fee12344fee12334fff00000fff00000fde11205fde01205ffe00105fff00104fff00016ffe00136fff00001fff00001;
assign testcases[629] = 512'hfde11344fde13344ffd01344ffd01344fdd13344fdd13434fff00000fff00000fde11305fde11305ffd00105fff00104fff00117fed00247fff00001fef00001;
assign testcases[630] = 512'hfde11454fde13454ffc01445ffd01345fdd13455fdd13445fff00000fff00001fdd11306fdd11306ffc00106fff00105ffe00117fec01257fff00001fef00001;
assign testcases[631] = 512'hfcd21454fcd14464ffc01455ffc01455fdc14465fdc14555fff00000fff00001fcd11306fcd12306ffc00106fff00105ffe00128fec01267fff00001fef00001;
assign testcases[632] = 512'hfcd21565fcd14465ffb01455ffc01465fcc14576fcc24556fff00000fff00001fcc12406fcc12406ffb01106fff01105ffe00128feb01368fff00001fef00001;
assign testcases[633] = 512'hfcd21575fcd14575ffb01566ffb01466fcb14576fcb25666fff00000fff00001fcc12407fcc12407ffb01107fff01106ffe00128feb01378fff00001fef00001;
assign testcases[634] = 512'hfbc21575fcc25575fea02566feb02576fcb15686fcb25667fff00001fff00001fcc12407fcc12507ffa01107ffe01106ffd00129fda01379fff00001fef00001;
assign testcases[635] = 512'hfbc21675fbc25686fea02577fea02576fbb15687fbb26777fff00001fff00001fbb12507fbb12507fea01108ffe01107ffd00129fda01389fff00001fef00001;
assign testcases[636] = 512'hfbc31686fbc25686fe902577fea02577fba15697fba26777fff00001fff00001fbb12508fbb12507fea01108ffe01107ffd00129fd901399fff00001fef00001;
assign testcases[637] = 512'hfbc21696fbb25696fe901687fea01587fba157a7fba26787fff12201fff12211fbb12508fbb12508fe901208ffe01107ffd00139fd901399fff01201fef01101;
assign testcases[638] = 512'hfef00112fef00112fff00112fff00112fff00112fff00112fff00000fff00000fef00004fef00103fff00003fff00002fff00005fff00014fff00001fff00000;
assign testcases[639] = 512'hfef00122fef01122fff00122fff00122fef01123fef01123fff00000fff00000fef00104fef00104fff00003fff00003fff00015fff00125fff00001fff00000;
assign testcases[640] = 512'hfef00132fef01132ffe00223fff00133fef01133fef01223fff00000fff00000fef00104fef00104fff00004fff00003fff00015fff00135fff00001fff00001;
assign testcases[641] = 512'hfdf10233fdf01233ffe01233ffe01233fef01233fef11233fff00000fff00000fef01104fef01104ffe00104fff00103fff00016ffe00135fff00001fff00001;
assign testcases[642] = 512'hfdf10233fdf12243ffe01233ffe01233fee02244fee12234fff00000fff00000fde01205fde01205ffe00104fff00104fff00016ffe00146fff00001fef00001;
assign testcases[643] = 512'hfde11343fde12343ffd01344ffd01344fde12344fde12344fff00000fff00000fde11205fde01205ffd00105fff00104fff00017fed00246fff00001fef00001;
assign testcases[644] = 512'hfde11354fde13354ffc01344ffd01354fdd13455fdd13445fff00000fff00001fdd11306fdd11305ffd00105fff00105fff00117fed00257fff00001fef00001;
assign testcases[645] = 512'hfcd21464fcd13464ffc01455ffc01355fdd13465fdd14455fff00000fff00001fcd11306fcd11306ffc00106fff00105ffe00127fec01267fff00001fef00001;
assign testcases[646] = 512'hfcd21465fcd14465ffb01455ffc01465fcc14575fcc24555fff00000fff00001fcd12306fcd12406ffb01106fff01105ffe00128feb01268fff00001fef00001;
assign testcases[647] = 512'hfcd21575fcd14575ffb01566ffb01466fcc14576fcc25666fff00000fff00001fcc12407fcc12407ffb01107fff01106ffe00128feb01378fff00001fef00001;
assign testcases[648] = 512'hfbc21575fcc15575fea01566feb01476fcb15686fcb25666fff00001fff00001fcc12407fcc12407ffa01107ffe01106ffd00129fda01388fff00001fef00001;
assign testcases[649] = 512'hfbc21686fbc25586fea02577fea01577fbb15697fbb25777fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fda01389fff00001fef00001;
assign testcases[650] = 512'hfbc32686fbc25686fe902677fea02577fba15797fba26777fff00001fff00001fbb22508fbb12508fe901108ffe01107ffd0012afd901399fff00001fef00001;
assign testcases[651] = 512'hfbb31686fbb25696fe902687fe902687fba157a8fba26787fff11201fff12211fbb12508fbb12508fe901208ffe01207ffd0013afd80149afff01201fef01101;
assign testcases[652] = 512'hfbc215a5fbc155a5fe902677fea02586fbb145b7fbb25687fff01101fff01111fbb12407fbb12407fea01108ffe01106ffd00139fda013a9fff01101fef01101;
assign testcases[653] = 512'hfbc21586fbc25596fe901577fea01587fba14697fbb25677fff00001fff00101fbb12407fbb12507fea01108ffe01107ffd00129fd901399fff00001fef00001;
assign testcases[654] = 512'hfbc21585fbc25585fe902577fea01576fbb15697fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01106ffd00129fda01399fff00001fef00001;
assign testcases[655] = 512'hfef00012fef00012fff00012fff00012fff00012fff00012fff00112fff01112fef00003fef00003fff00003fff00002fff00005fff00014fff00103fef00102;
assign testcases[656] = 512'hfef00012fef00012fff00112fff00112fff00012fff00012fef01113fff01113fef00003fef00003fff00003fff00003fff00005fff00014ffe01103fef01103;
assign testcases[657] = 512'hfef00012fef00012fff00123fff00123fff00012fff00012fee11113fee11114fef00004fef00004fff00004fff00003fff00005fff00014fee01104fde01104;
assign testcases[658] = 512'hfef00012fef00012fff00123fff00123fff00013fef00013fdd11214fed12215fef00004fef00004fff00004fff00003fff00005fff00015fed01205fdd01204;
assign testcases[659] = 512'hfef00012fef00012ffe00123fff00123fef00023fef00013edd12215fdc12215fef00004fef00004fff00004fff00003fff00005fff00025fec01306edd12205;
assign testcases[660] = 512'hfef00123fef00123ffe00124ffe00124fef00123fef00113ecc12315fdc12316fef00004fef00004ffe00005fff00004fff00005fff00025fdb01306ecc12306;
assign testcases[661] = 512'hfef00123fef00123ffe00134ffe00134fef00123fef00123ecc23316fdb13416fef00104fef00104ffe00005fff00004fff00015fff00025fdb02407ecc13406;
assign testcases[662] = 512'hfbbf2815fabf9815fe713926fe813826fa9f9a17fa9faa17fff00000fff00000fbab4707fba84707fe701207ffe01206fff14206fff00a04fff00001feff9201;
assign testcases[663] = 512'hfef32712fef27712ffe02723fff02623fef27813fef38913fff00000fff00000fef23604fef23604fff01204fff01203fcc27404fadfec04fff00001fff86100;
assign testcases[664] = 512'hfbb32787fbb27787fe802778fe902688fb927898fb938878fff00000fff00001fba23609fba23608fd801209ffe01208eee27457fff00a04fdf00001ecf00001;
assign testcases[665] = 512'h25b3277758b2778700002778002026780092789805938978def00000fff0000147a2360906a23608000012098bb01208fee14225f0800a19ccf00001bbf00001;
assign testcases[666] = 512'hfaa8fe98faa9fa98fe6afe8afe7aff9afa84dbaafa88fc8afff11101fff11101fa9f6afafa9f7bfafe7fc7fcffdfe8fb37b385fcfc60fc2afff01231fef011f1;
assign testcases[667] = 512'hfaa32737faa27737fc602759fb714859fa84ba39fa88db29fff00000fff01100fa986a09fa956a099471340a000134090004841cfc64273bc5d00101c9f00001;
assign testcases[668] = 512'hf9b84a25fbc5c925fe814b36feb13b25fde3dd14fde5dd14fff00000fff00000fef66903fef11103fff01103fff12302fff12204fff01114fff01100fff01000;
assign testcases[669] = 512'hfef84e13fef6fd13ffe14e13ffe14d14fef4de13fef6ef13fff00000fff01100fef46a05fef36b04fff12304fff12404fff00004fff02715fff00101fff00000;
assign testcases[670] = 512'hfef00001fef00001fff00001fff00001fff00002fff00002fff00000fff00000fef00003fef00003fff00002fff00001fff00004fff00004fff00000fff00000;
assign testcases[671] = 512'hfef00001fef00001fff00001fff00001fff00002fff00002fff00000fff00000fef00003fef00003fff00002fff00001fff00004fff00004fff00000fff00000;
assign testcases[672] = 512'hfef00001fef00001fff00001fff00001fff00002fff00002fff00000fff00000fef00003fef00003fff00002fff00001fff00004fff00004fff00000fff00000;
assign testcases[673] = 512'hfef00001fef00001fff00001fff00001fff00002fff00002fff00000fff00000fef00003fef00003fff00002fff00001fff00004fff00004fff00000fff00000;
assign testcases[674] = 512'hfef00001fef00001fff00001fff00001fff00002fff00002fff00000fff00000fef00003fef00003fff00002fff00001fff00004fff00004fff00000fff00000;
assign testcases[675] = 512'hfef00001fef00001fff00001fff00001fff00002fff00002fff00000fff00000fef00003fef00003fff00002fff00001fff00004fff00004fff00000fff00000;
assign testcases[676] = 512'hfef00001fef00001fff00001fff00001fff00002fff00002fff00000fff00000fef00003fef00003fff00002fff00001fff00004fff00004fff00000fff00000;
assign testcases[677] = 512'hfef00001fef00001fff00001fff00001fff00002fff00002fff00000fff00000fef00003fef00003fff00002fff00001fff00004fff00004fff00000fff00000;
assign testcases[678] = 512'hfef10112fef01112ffe01323ffe01323fff01112fef01112fef01111fff01111fef01104fef01103fff00103fff01103fff00005fff00014fff00101fef01101;
assign testcases[679] = 512'hfef10112fef01112ffe01323ffe01323fef01112fef01112fff01111fff01111fef00104fef00104fff00104fff00103fff00005fff00014fff00101fef01101;
assign testcases[680] = 512'hfef10123fef01122ffd01434ffe01434fef01123fef01113fef11112fff01112fef01104fef01104ffe00104fff01104fff00005fff00125fff01102fef01102;
assign testcases[681] = 512'hfef10223fef01223ffd01435ffd01445fef01223fef11223fee12222fee12212fef01104fef01104ffe00105fff01105fff00015fff00125ffe01202fef01102;
assign testcases[682] = 512'hfdf10223fdf12223ffc01545ffc01545fef02223fef12223fde12223fee12222fef01104fef01104ffd00105fff01105fff00016fff00125fee01202fde02202;
assign testcases[683] = 512'hfde11233fde12233ffb02546ffc02556fee02234fee12224fdd12323fed12223fde11105fee01205ffd01106fff01106fff00016ffe00125fee01203fde02202;
assign testcases[684] = 512'hfde11334fde12344ffa02657ffb02657fde12234fde12334fdd23334fdd13323fde11205fde01205ffc01107ffe01207fff00016ffe00136fed02303fdd13303;
assign testcases[685] = 512'hfcd11344fde13344fe902768fea02768fdd12345fdd13334ecc24434fdc24434fde11206fde11205ffb01107ffe01207fff00016ffd00136fec02304fcd13304;
assign testcases[686] = 512'hfcd11445fcd13455fe802868fe902778fdd13345fdd13335ecb35535fdb24534fdd11206fdd11306ffa01108ffe01208fff00017fed00146fec02404fcc14404;
assign testcases[687] = 512'hfcd21455fcd13455fe803979fe802879fdc13455fdd13445ebb35535fdb25535fcd11306fcd11306fea01208ffe01209fff00017fed00247fdb03405ecc14404;
assign testcases[688] = 512'hfbc21556fcc13455fe71397afe81388afcc13456fcc13446eba36636fcb26535fcc11307fcc11307fe901209ffe0120affe00017fec00247fdb03505ecb15505;
assign testcases[689] = 512'hfbc21566fbc14566fe613a8afe71398afcc14466fcc13546eba46636fca36646fcc11307fcc11307fe80120affd0120affe00118fec00257fdb13505ebb15505;
assign testcases[690] = 512'hfbb21566fbb14566fe513a8bfe71399bfcb14566fcb14556eba47746fca37646fcc11307fcc12407fe80120affd0120bffe00118feb00258fda13606ebb16605;
assign testcases[691] = 512'hfab21667fbb14577fe513a8bfe61399bfcb14567fcb24557ea947747fc937746fcb11408fbb12407fe70120affd0130bffe00118feb01268fda14606eba26606;
assign testcases[692] = 512'hfef00112fef01112ffe01323ffe01323fff01112fef01112fff01111fff01111fef00104fef00104fff00104fff00103fff00005fff00014fff00101fef01101;
assign testcases[693] = 512'hfef10123fef01122ffd01434ffe01334fef01123fef01113fef11112fff01112fef00104fef00104ffe00104fff00104fff00005fff00125fff01102fef01102;
assign testcases[694] = 512'hfef10223fef01223ffd01435ffd01445fef01123fef11223fee12212fee11212fef01104fef01104ffe00105fff01105fff00015fff00125ffe01202fef01102;
assign testcases[695] = 512'hfdf10233fdf01233ffc01545ffc01445fef01223fef11223fde12223fee12222fef01105fef01104ffd00105fff01105fff00016fff00125fee01202fde02202;
assign testcases[696] = 512'hfde11233fde12233ffb01546ffc01556fee02234fee12224fdd12323fed12223fde01105fde01205ffd00106fff01106fff00016ffe00125fee01203fde02203;
assign testcases[697] = 512'hfde11344fde12344ffa02657ffb02657fee12234fee12334edc23324fdd13323fde11205fde01205ffc01107fff01207fff00016ffe00136fed02303fdd13303;
assign testcases[698] = 512'hfcd11344fde12344fe902768fea02768fdd12345fdd12335ecc24434fdc24434fde11206fde11206ffb01107ffe01208fff00017ffe00136fec02304fcd13304;
assign testcases[699] = 512'hfcd11455fcd13455fe802868fe902778fdd13345fdd13335ecb35535fdb24534fdd11206fdd11306ffa01208ffe01208fff00017fed00146fec02404ecc14404;
assign testcases[700] = 512'hfcd21455fcd13455fe803979fe902879fdd13455fdd13445ebb35535fdb25535fcd11306fcd11306ffa01209ffe01209fff00017fed00247fdb03405ecc14404;
assign testcases[701] = 512'hfbc21556fcc13455fe71397afe80388afcc13456fcc13446eba36636fcb26535fcc11307fcc11307fe901209ffe0120affe00017fec00247fdb03505ecb15505;
assign testcases[702] = 512'hfbc21566fbc14566fe613a8afe71398afcc14456fcc14546eba46646fca36646fcc11307fcc12407fe90120affd0120affe00118fec00257fdb13505ebb15505;
assign testcases[703] = 512'hfbb21666fbb14566fe513a8bfe71399bfcb14566fcb14556eba47746fca37646fcc11407fcc12407fe80120affd0120bffe00118feb01258fda13606ebb16605;
assign testcases[704] = 512'hfbb21667fbb14677fe513b8bfe61399bfcb14567fcb24557ea947747fc937746fbb12408fbb12408fe70120bffd0130bffe00118feb01258fda14606eba26606;
assign testcases[705] = 512'hfef00112fef01112ffe01223ffe01223fef01112fef01112fff01111fff00111fef00104fef00104fff00004fff00103fff00005fff00014fff00101fef00001;
assign testcases[706] = 512'hfef00123fef01122ffd01334ffe01334fef01123fef01113fef11112fff01112fef00104fef00104ffe00104fff00104fff00005fff00025fff01102fef01102;
assign testcases[707] = 512'hfef10223fef01223ffc01435ffd01445fef01123fef01223fee12222fee11222fef00104fef01104ffd00105fff00105fff00015fff00125ffe01102fef01102;
assign testcases[708] = 512'hfdf10223fdf01223ffc01545ffc01445fef01223fef11223fde12223fee12222fef01105fef01104ffd00105fff01105fff00016fff00125fee01202fde02202;
assign testcases[709] = 512'hfde11233fde02233ffb01546ffc01556fee02234fee12224fdd12323fed12223fde01105fde01205ffd00106fff01106fff00016ffe00125fee01203fde02203;
assign testcases[710] = 512'hfde11334fde12334ffa02757ffb02657fee12234fee12334fdc23324fdd13323fde11205fde01205ffc01107ffe01207fff00016ffe00136fed02303fdd13303;
assign testcases[711] = 512'hfcd11344fdd13344fe902768fea02768fdd12345fdd13335ecc24434fdc24434fdd11206fdd11206ffb01107ffe01208fff00017fed00136fec02304fcd13304;
assign testcases[712] = 512'hfcd11445fcd13455fe802869fe902778fdd13345fdd13435ecb35535fdb24534fdd11306fdd11306ffa01208ffe01208fff00017fed00147fec02404fcc14404;
assign testcases[713] = 512'hfcc21555fcd13455fe803979fe803879fdc13455fdc13445ebb35545fdb25535fcd11306fcd11306ffa01209ffe01209ffe00017fec00247fdb03405ecc14404;
assign testcases[714] = 512'hfbc21556fcc14556fe71397afe81388afcc13456fcc14446eba36646fca26645fcc11307fcc11307fe901209ffd0120affe00118fec00247fdb03505ecb15505;
assign testcases[715] = 512'hfbc21566fbc14566fe613a8afe71398afcc14456fcc14546eba46646fca36646fcc11307fcc12407fe80120affd0120affe00118fec00258fdb13505ebb15505;
assign testcases[716] = 512'hfbb21667fbb14566fe513a8bfe61399bfcb14567fcb24557eba47746fca37646fbb12408fcb12408fe80120affd0130bffe00118feb01258fda13606ebb16505;
assign testcases[717] = 512'hfab21667fbb14677fe513b8cfe613a9bfbb14567fbb24657ea947747fc937746fbb12408fbb12408fe70120bffd0130bffe00118feb01268fda14606ebb26606;
assign testcases[718] = 512'hfef00112fef01112ffe01323ffe01323fef01112fef01112fff01111fff01111fef00104fef00104fff00104fff00103fff00005fff00014fff00101fef00101;
assign testcases[719] = 512'hfef10123fef01122ffd01434ffd01334fef01123fef01113fef11112fff01112fef01104fef01104ffe00104fff01104fff00005fff00125fff01102fef01102;
assign testcases[720] = 512'hfdf10223fef01223ffc01535ffd01445fef01223fef11223fee12222fee11222fef01104fef01104ffd00105fff01105fff00015fff00125ffe01102fef01102;
assign testcases[721] = 512'hfdf10233fdf12233ffc01546ffc01545fef02223fef12223fde12223fee12222fef01105fef01205ffd00105fff01105fff00016fff00125fee01202fde02202;
assign testcases[722] = 512'hfde11233fde12233ffb02646ffc02556fee12234fee12224fdd12323fed12223fde11205fde01205ffc01106fff01106fff00016ffe00125fee01203fde02202;
assign testcases[723] = 512'hfde11344fde12344ffa02757ffb02667fde12334fde12334fdd23334fdd13333fde11205fde11205ffb01107ffe01207fff00016ffe00136fed02303fdd13303;
assign testcases[724] = 512'hfcd11445fdd13344fe902868fea02768fdd13345fdd13335ecc24434fdc24434fdd11206fdd11306ffb01108ffe01208fff00017fed00136fec02304fcd13304;
assign testcases[725] = 512'hfcd21455fcd13455fe802869fe902879fdd13445fdd13435ecb35545fdb24434fcd11306fcd11306ffa01208ffe01209fff00017fed00247fec02404fcc14404;
assign testcases[726] = 512'hfcc21555fcc13455fe703979fe813879fdc13456fcc13446ecb35545fdb25535fcc11307fcc11307fe901209ffe01209ffe00017fec00247fdb03405ecc14404;
assign testcases[727] = 512'hfbc21556fcc14556fe613a7afe71398afcc14456fcc14546eba36645fcb26545fcc11307fcc12407fe901209ffd0120affe00118fec00247fdb03505ecc15505;
assign testcases[728] = 512'hfbb21666fbc14566fe613a8bfe71398bfcb14556fcb24546eba46646fca36646fcc12407fcc12407fe80120affd0130affe00118feb01258fdb13505ebb15505;
assign testcases[729] = 512'hfbb21667fbb14666fe513a8bfe61399bfcb14567fcb24557eba47746fca37646fbb12408fbb12408fe80120affd0130bffe00118feb01258fda13606ebb16505;
assign testcases[730] = 512'hfab21667fbb15677fe413b8cfe513a9cfba14567fbb24657ea947746fc937746fbb12408fbb12408fe70120bffd0130cffe00119fea01258fda14606ebb16606;
assign testcases[731] = 512'hfef00112fef01112ffe01323ffe01223fef01113fef01112fff01111fff00111fef00104fef00104fff00104fff00103fff00005fff00014fff00101fef00001;
assign testcases[732] = 512'hfef10223fef01122ffd01434ffd01334fef01123fef01113fef11112fff01112fef00104fef01104ffe00104fff00104fff00005fff00115fff01102fef01102;
assign testcases[733] = 512'hfef10223fef01223ffd01435ffd01445fef01223fef11213fee12222fee11222fef01104fef01104ffd00105fff01105fff00005fff00125ffe01102fef01102;
assign testcases[734] = 512'hfdf10223fdf12223ffc01545ffc01445fef02223fef12223fde22223fee12222fef01105fef01204ffd00105fff01105fff00016fff00125fee01202fde02202;
assign testcases[735] = 512'hfde11233fde12233ffb02546ffc02556fee02224fee12224fdd12323fed12223fde11205fde01205ffd01106fff01106fff00016ffe00125fee01203fde02202;
assign testcases[736] = 512'hfde11334fde12334ffa02657ffb02657fee12234fee12324edc23324fdd13323fde11205fde01205ffc01106fff01207fff00016ffe00136fed02303fdd13303;
assign testcases[737] = 512'hfcd11344fde13344fe902768fea02767fdd12334fdd13334ecc24424fdc24424fde11206fde11206ffb01107ffe01207fff00017ffd00136fec02304fcd13304;
assign testcases[738] = 512'hfcd11445fcd13445fe902868fe902778fdd13345fdd13335ecb35535fdb24524fdd11206fdd11306ffa01108ffe01208fff00017fed00147fec02404fcc14404;
assign testcases[739] = 512'hfcd21455fcd13455fe802879fe902879fdd13445fdd13445ebb35535fdb25525fcd11306fcd11306ffa01208ffe01209fff00017fed00247fdb03405ecc14404;
assign testcases[740] = 512'hfbc21556fcc13455fe70397afe80388afcc13456fcc13446eba36636fca26535fcc11307fcc11307fe901209ffe0120affe00118fec00247fdb03505ecb15505;
assign testcases[741] = 512'hfbc21556fbc14556fe61397afe71398afcc14456fcc14546eba46636fca36636fcc11307fcc12407fe80120affd0120affe00118fec00258fdb13505ebb15505;
assign testcases[742] = 512'hfbb21666fbb14566fe613a8bfe71398bfcb14556fcb24546eba47736fca37636fcb12407fcb12407fe80120affd0130bffe00118feb01258fda13506ebb16505;
assign testcases[743] = 512'hfbb21667fbb14667fe513a8bfe61399bfcb14567fcb24557ea947737fc937736fbb12408fbb12408fe70120bffd0130bffe00118feb01258fda14606eba26606;
assign testcases[744] = 512'hfbc21586fbc25586fe901577fea01577fba15697fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fda01389fff00001fef00001;
assign testcases[745] = 512'hfbc21586fbc25585fe901577fea01587fba15697fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fd901399fff00001fef00001;
assign testcases[746] = 512'hfbc21686fbc25585fe901577fea01576fba15697fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fd901389fff00001fef00001;
assign testcases[747] = 512'hfbc21586fbc25585fe901577fea01576fba15697fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fd901399fff00001fef00001;
assign testcases[748] = 512'hfbc21675fbc25685fe902577fea02576fba15687fbb25677fff00001fff00001fbb12507fbb12507fea01108ffe01106ffd00129fda01389fff00001fef00001;
assign testcases[749] = 512'hfbc21585fbc15595fea01576fea01476fbb14696fcb25676fff00001fff00001fbb12407fbb12407fea01107ffe01106ffd00129fda01398fff00001fef00001;
assign testcases[750] = 512'hfbc21586fbc14596fe901577fea01487fba146a7fbb25677fff00001fff00001fbb12407fbb12407fea01108ffe01107ffd00129fda01399fff00001fef00001;
assign testcases[751] = 512'hfbc32635fbc26635fe902636fea02546fba26646fbb26736fff00001fff00001fbb22507fbb13507fea01207ffe01206ffd00119fd901338fff00001fef00001;
assign testcases[752] = 512'hfbc21675fbc25585fe902577fea01577fba15687fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fd901389fff00001fef00001;
assign testcases[753] = 512'hfbc21565fbc25565fe902566fea01576fba15677fbb25666fff00001fff00001fbb12407fbb12507fea01107ffe01106ffd00129fda01379fff00001fef00001;
assign testcases[754] = 512'hfbc21555fbc15565fea01566fea01576fbb15666fbb25656fff00001fff00001fbb12407fbb12507fea01107ffe01106ffd00129fda01369fff00001fef00001;
assign testcases[755] = 512'hfbc21585fbc25595fe901577fea01586fba15697fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fda01399fff00001fef00001;
assign testcases[756] = 512'hfbc21686fbc25586fe902577fea01587fba15697fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fd901399fff00001fef00001;
assign testcases[757] = 512'hfbc21686fbc25596fe902577fea01587fba15697fbb25677fff00001fff00001fbb12407fbb12507fea01108ffe01107ffd00129fd901399fff00001fef00001;
assign testcases[758] = 512'hfbb32796fbb26696fe802787fe902687fba157a7fba26887fff12201fff12311fbb22508fbb12608fe901208ffe01207ffd0013afd8014a9fff01201fef02201;
assign testcases[759] = 512'hfbb21696fbb25696fe902687fe902587fba157a7fba26787fff01101fff01111fbb12508fbb12508fe901208ffe01107ffd0013afd9014a9fff01101fef01101;
assign testcases[760] = 512'hfbc215a5fbc145b5fea01586fea01586fcb146b6fcb25696fff00001fff00001fbc12407fcc12407fea01107ffe01106ffd00139fda013b8fff00001fef00001;
assign testcases[761] = 512'hfbc21585fbc14595fea01576fea01486fbb14596fbb24676fff00001fff00001fbb12407fcc12407fea01107ffe01106ffd00129fda01398fff00001fef00001;
assign testcases[762] = 512'hfbc21565fbc25565fe901566fea01576fba15677fbb25656fff00000fff00001fbb12407fbb12407fea01107ffe01106ffd00129fda01368fff00001fef00001;
assign testcases[763] = 512'hfbc21586fbc15585fe901577fea01586fba15697fbb25677fff00000fff00001fbb12407fbb12407fea01108ffe01107ffd00129fda01389fff00001fef00001;
assign testcases[764] = 512'hfbc21696fbc25596fe901577fea02587fba156a7fba25687fff00001fff00001fbb12408fbb12507fe901108ffe01107ffd00139fd901399fff00001fef00001;
assign testcases[765] = 512'hfbb21676fbb25686fe902677fea02577fba15687fba26777fff00000fff00001fbb12508fbb12508fe901108ffe01107ffd00129fd901389fff00001fef00001;
assign testcases[766] = 512'hfab32797fab27797fe802788fe802688fa9268a8fa937988fff01101fff01111faa23609fba13609fe801209ffe01208ffc0113bfd70149afff00101fef00101;
assign testcases[767] = 512'hfef00112fef01112fff00112fff00112fef01113fef01112fff00000fff00000fef00104fef00104fff00003fff00002fff00005fff00015fff00001fff00000;
assign testcases[768] = 512'hfef00123fef01122ffe00223fff00223fef01123fef01223fff00000fff00000fef00104fef00104fff00004fff00003fff00016fff00125fff00001fff00000;
assign testcases[769] = 512'hfdf10233fdf01233ffe01233ffe01233fee02234fee12224fff00000fff00000fdf01205fef01205ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[770] = 512'hfde11233fde12233ffd01334ffe01234fee12334fee12334fff00000fff00000fde11205fde01205ffd00105fff00104fff00016ffe00136fff00001fff00001;
assign testcases[771] = 512'hfde11334fde12333ffd01334ffd01334fde12344fde12334fff00000fff00000fde11205fde01205ffd00105fff00104fff00017fed00236fff00001fff00001;
assign testcases[772] = 512'hfde11444fde13444ffc01445ffc01445fdd13445fdd14445fff00000fff00000fdd11306fdd11306ffc00106fff00105ffe00117fec01247fff00001fef00001;
assign testcases[773] = 512'hfcd21555fcd14455ffb01546ffc01455fcc14556fcc24546fff00000fff00000fcd12407fcd12406ffb01107fff01106ffe00118feb01358fff00001fef00001;
assign testcases[774] = 512'hfcd21555fcd25555fea02556ffb02556fcb15666fcb25656fff00000fff00000fcc12407fcc12407ffb01107fff01106ffe00129feb01358fff00001fef00001;
assign testcases[775] = 512'hfbc31666fcc26666fea02657fea02567fcb15667fcb26757fff00000fff00001fcc22507fcc12507fea01208ffe01207ffd00129fda01369fff00001fef00001;
assign testcases[776] = 512'hfbc32666fbc26666fe902667fea02667fba26777fba37757fff00000fff00001fbb22508fbb13508fe901208ffe01207ffd0012afd901469fff00001fef00001;
assign testcases[777] = 512'hfbb32776fbb27776fe802768fe902678fba26888fba37868fff00000fff00001fba23508fbb13608fe901209ffe01208ffd0112afd80147afff00001fef00001;
assign testcases[778] = 512'hfbb32777fbb27777fe802778fe902678fb927888fa938968fff00000fff00001fba23609fba23609fe801209ffe01208ffd0112bfd80148bfff00001fef00001;
assign testcases[779] = 512'hfab42877fab38887fe702879fe802778fa827989fa938979fff00000fff00001fba23609fba23709fe70120affe01209ffc0112bfd70158bfff00001fef00001;
assign testcases[780] = 512'hfef00112fef01112fff00123fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00005fff00115fff00001fff00000;
assign testcases[781] = 512'hfef10223fef01223ffe01223ffe01223fef01223fef11223fff00000fff00000fef01104fef01104ffe00104fff00103fff00016ffe00125fff00001fff00000;
assign testcases[782] = 512'hfdf10233fdf12233ffe01334ffe01234fee12234fee12324fff00000fff00000fde11205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[783] = 512'hfde11333fde12333ffd01334ffd01334fee12334fde12334fff00000fff00000fde11205fde01205ffd00105fff00104fff00017ffd00236fff00001fff00001;
assign testcases[784] = 512'hfde11334fde13334ffd01434ffd01334fdd13344fdd13435fff00000fff00000fde11306fde11305ffd00105fff00105fff00117fed00237fff00001fff00001;
assign testcases[785] = 512'hfcd21444fdd14444ffc01445ffc01445fdd13445fdd14545fff00000fff00000fdd11306fdd12306ffc01106fff00105ffe00118fec01247fff00001fef00001;
assign testcases[786] = 512'hfcd21555fcd14555ffb01546ffc01456fcc14556fcc25646fff00000fff00000fcc12407fcc12407ffb01107fff01106ffe00118feb01358fff00001fef00001;
assign testcases[787] = 512'hfcc21555fcc25555fea02556feb02556fcb15666fcb25656fff00000fff00000fcc12407fcc12507ffa01107ffe01106ffe00129fea01369fff00001fef00001;
assign testcases[788] = 512'hfbc32666fbc26666fea02657fea02567fcb15667fbb26757fff00000fff00001fcb22508fcb12507fea01208ffe01107ffd00129fda01369fff00001fef00001;
assign testcases[789] = 512'hfbc32666fbc26666fe902667fea02667fba26777fba37857fff00000fff00001fbb23508fbb13508fe901208ffe01207ffd0012afd90147afff00001fef00001;
assign testcases[790] = 512'hfbb32766fbb27776fe802768fe902668fb927878fba37868fff00000fff00001fba23608fbb13608fe901209ffe01208ffd0112afd80147afff00001fef00001;
assign testcases[791] = 512'hfbb32777fbb27777fe802778fe902678fb927888fa938968fff00000fff00001fba23609fba23609fe801209ffe01208ffc0112bfd80147bfff00001fef00001;
assign testcases[792] = 512'hfab42877fab38787fe702779fe802778fa827989fa938979fff00000fff00001faa23609faa23609fe80120affe01209ffc0112bfd70158bfff00001fef00001;
assign testcases[793] = 512'hfef00112fef01112fff00213fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00005fff00115fff00001fff00000;
assign testcases[794] = 512'hfef10223fef01223ffe01223ffe01223fef01223fef11223fff00000fff00000fef01104fef01204ffe00104fff00103fff00016ffe00125fff00001fff00000;
assign testcases[795] = 512'hfdf10233fdf12233ffe01334ffe01233fee12234fee12324fff00000fff00000fde01205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[796] = 512'hfde11333fde12333ffd01334ffd01334fde12334fde12334fff00000fff00000fde11205fde01205ffd00105fff00104fff00017fed00236fff00001fff00001;
assign testcases[797] = 512'hfde11334fde13334ffd01434ffd01334fdd13344fdd13434fff00000fff00000fde11305fde11305ffd00105fff00104fff00117fed00237fff00001fff00001;
assign testcases[798] = 512'hfdd21444fdd14444ffc01445ffc01445fdd14445fdd14545fff00000fff00000fdd11306fdd12306ffc01106fff01105ffe00118fec01247fff00001fef00001;
assign testcases[799] = 512'hfcd21555fcd14555ffb01546ffc01455fcc14556fcc25646fff00000fff00000fcc12407fcd12406ffb01107fff01106ffe00118feb01358fff00001fef00001;
assign testcases[800] = 512'hfcd21555fcd25555ffa02556ffb02556fcb15666fcb25656fff00000fff00000fcc12407fcc12507ffb01107fff01106ffe00129fea01369fff00001fef00001;
assign testcases[801] = 512'hfbc32666fcc26666fea02657fea02567fcb15667fcb26757fff00000fff00001fcb22508fcb12507fea01208ffe01107ffd00129fda01369fff00001fef00001;
assign testcases[802] = 512'hfbc32666fbc26666fe902667fea02667fba26777fba37857fff00000fff00001fbb23508fbb13508fe901208ffe01207ffd0012afd90147afff00001fef00001;
assign testcases[803] = 512'hfbb32766fbb27776fe802768fe902678fba26878fba37868fff00000fff00001fbb23508fbb13608fe901209ffe01208ffd0112afd80147afff00001fef00001;
assign testcases[804] = 512'hfbb32777fbb27777fe802768fe902678fb927888fb938968fff00000fff00001fba23609fba23608fe801209ffe01208ffd0112bfd80147afff00001fef00001;
assign testcases[805] = 512'hfab42777fab38777fe702779fe802778fa927889fa938979fff00000fff00001faa23609faa23609fe80120affe01208ffc0112bfd70158bfff00001fef00001;
assign testcases[806] = 512'hfef00112fef01112fff00112fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00005fff00115fff00001fff00000;
assign testcases[807] = 512'hfef10223fef01223ffe01223ffe01223fef01223fef11223fff00000fff00000fef01104fef01204ffe00104fff00103fff00016fff00125fff00001fff00000;
assign testcases[808] = 512'hfdf10223fdf12223ffe01324ffe01233fee12234fee12324fff00000fff00000fde11205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[809] = 512'hfde11333fde12333ffd01334ffd01334fde12334fde12324fff00000fff00000fde11205fde01205ffd00105fff00104fff00017fed00236fff00001fff00001;
assign testcases[810] = 512'hfde11334fde13334ffd01334ffd01334fdd13334fdd13435fff00000fff00100fde11305fde11305ffd00105fff00104fff00117fed00237fff00101fff00001;
assign testcases[811] = 512'hfcd21444fcd14444ffc01445ffc01445fdd14445fdd14545fff00000fff00000fcd11306fdd12306ffc01106fff01105ffe00118fec01247fff00001fef00001;
assign testcases[812] = 512'hfaa42987faa39988fe613a79fe713989fa829b99fa84ab7afff54301fff54411fa9dff0afa9aff09fe66ff0bffd5ff09ffc0442bfc61af8cfff13401fef14300;
assign testcases[813] = 512'hfab42867fab38867fe702869fe802778fa828979fa938969fff00000fff00001fba23609fba23609fe70120affe01209ffd0112afd70157bfff00001fef00001;
assign testcases[814] = 512'hfab42877fab38877fe702879fe802778fa828989fa939969fff00000fff00001faa23609fba23709fe70120affe01209ffd0112afd70158bfff00001fef00001;
assign testcases[815] = 512'hfab42877fab38877fe702879fe802778fa828989ea939969fff00000fff00001faa23609eaa23709fe70120affe01209ffc0112bfc70158bfff00001fef00001;
assign testcases[816] = 512'hfaa42987faa39988fe602979fe712889fa828a99fa84ab79fff11111fff11211fa92470afa924709fe60120bffd01209ffc0112bfc60159cfff01201fef02201;
assign testcases[817] = 512'hfaa42867faa39867fe602879fe702779fa728a79f9849a59fff00001fff01101fa92370afa924709fe60120bffd012096530112bfc60156cfff01101f5e01101;
assign testcases[818] = 512'hfab42877fab38877fe702879fe802779fa828989fa939969fff00000fff00001faa23609fba23709fe70120affe01209ffd01129fd70157bfff00001fef00001;
assign testcases[819] = 512'heab42867eab38867fe712879fe812778e9828979d9939969fff00000fff00001eaa23609daa23709fe70120affe01209ffd01129dc70157bfff00001fef00001;
assign testcases[820] = 512'hfab42877fab38877fe702879fe802779fa828989fa939969fff00000fff00001faa23609fba23709fe70120affe01209ffd0113afd70158bfff00001fef00001;
assign testcases[821] = 512'hfab42877fab38877fe702879fe802779fa828989fa939969fff00000fff00001faa23609fba23709fe70120affe01209ffd0112afd70158bfff00001fef00001;
assign testcases[822] = 512'hfaa42988faa39988fe60297afe702889fa728a9afa84ab7afff11101fff11201fa92470afa92470afe60120bffd01209ffd0113afc60158cfff01201fef01101;
assign testcases[823] = 512'hfaa42878faa39888fe60297afe702889fa728a9af9849a7afff00101fff01101fa92470afa924709fe60120bffd012098860112af460158ce7d01101fef01101;
assign testcases[824] = 512'hfef42757fef38757fff02768fff02768fff37968fff48958fff00000fff00001fef33609fef23609fff01209fff01208ffffff25fffffb04fff00001fff00001;
assign testcases[825] = 512'hfab22515fbb26515fe7ffe26fe8ffe26fa925616fa945616fff00000fff00000fba42407fba32407fe8c7407ffea8506fff12104f6f00b04fff00001fef00000;
assign testcases[826] = 512'hfab42777fab38777fe702779fe802778fa927989fa938968fff00000fff00001fba23609fba23609fe80120affe01208fff00004fff00004fff00001fef00001;
assign testcases[827] = 512'hfab42777fbb38787fe702879fe802778fa927989fa938979fff00000fff00001fba23609fba23609fe80120affe01208fff00004fff00004fff00001fef00001;
assign testcases[828] = 512'hfaa42887faa38888fe602889fe702789fa828a99fa849a79fff11101fff11101fa92370afa924709fe70120bffd01209fff12136fff00004fff01201fef01101;
assign testcases[829] = 512'hfaa42887faa38887fe602879fe702789fa828a99fa849a79fff00001fff01101fa92370afa924709fe70120affd01209ffe01178fff00004fff00101fef01101;
assign testcases[830] = 512'hfaa42887faa38887fe602889fe702789fa828999fa839a79fff00001fff01101fa92370afa924709fe70120bffd01209eee11178fff00004fff00101fef00101;
assign testcases[831] = 512'hfaa42887faa38887fe602879fe702789fa828999fa849a79fff00001fff01101fa92370afa924709fe70120bffd01209ecd11157f2a00004fff00101fef00101;
assign testcases[832] = 512'hfbb32726fab27736fe802748fe802657fa927838fa937828fff00000fff00000fba23608fba13608fe801209ffe01208edf2430401800a04fffff301fef00001;
assign testcases[833] = 512'hfac32756fac27756fe802867fe902767fba26757eba37847fff12201fff13311fbb22507ebb12507fe901208ffe01208ffd00119eda01359fff02301fef13201;
assign testcases[834] = 512'hfbc32666fbb26666fe802778fe902677fba26777fba37867fff00001fff00101fbb22508fbb12507fe901208ffe01209ffd00129fd901379fff00101fef00001;
assign testcases[835] = 512'hfbc32676fbb26676fe802678fe902677fba26787fba37867fff00000fff00101fbb22508fbb12508fe901208ffe01209ffd00129fd901389fff00101fef00001;
assign testcases[836] = 512'hfbc32676fbb26676fe802678fe902677fba26788fba37878fff00000fff00001fbb22508fbb12508fe901208ffe01209ffd00129fd901389fff00101fef00001;
assign testcases[837] = 512'hfab32887fab27887fe702988fe802888fa927998fa938978fff24401fff24501fba23608fba13608fe801209ffd01309ffd0112afd80149afff03501fef14401;
assign testcases[838] = 512'hfab32777fab27777fe702778fe802688fa927888fa937868fff01101fff01101fba22508fba13608fe801209ffd01209ffd0012afd80147afff01101fef01101;
assign testcases[839] = 512'hfab32787fab27787fe702788fe802688fa927898fa937878fff01101fff01101fba23508fba13608fe801209ffd01209ffd0012afd80149afff01101fef01101;
assign testcases[840] = 512'hfab32787fab27787fe702788fe802688fa927898fa937878fff01101fff01101fba23508fba13608fe801209ffd01209ffd0012afd80149afff00101fef01101;
assign testcases[841] = 512'hfbb32656fbb26656fe802667fe902667fb926758fba26847fff00000fff00001fbb22508fbb12508fe901208ffe01208ffd0011afd901359fff00001fef00001;
assign testcases[842] = 512'hfbb32676fbb26676fe802678fe902677fb926788fba37868fff00000fff00001fbb22508fbb12508fe901208ffe01209ffd0012afd901489fff00001fef00001;
assign testcases[843] = 512'hfbb32676fbb26676fe802678fe902677fb926788fba37868fff00000fff00001fbb22508fbb12508fe901208ffe01209ffd0012afd901489fff00001fef00001;
assign testcases[844] = 512'hfbb32676fbb26676fe802678fe902677fb926888fba37868fff00000fff00001fbb22508fbb13508fe901208ffe01209ffd0012afd901489fff00001fef00001;
assign testcases[845] = 512'hfab32767fab27777fe702778fe802678fa927888fa937968fff11111fff11211fba23608fba13608fe901209ffd01209ffd0012afd80147afff01201fef01101;
assign testcases[846] = 512'hfab32757fab27757fe702778fe802678fa927868fa937858fff00001fff01101fba23508fba13608fe801209ffd01209ffc0012afd80146afff00101fef00101;
assign testcases[847] = 512'hfab32787fab27787fe702788fe802688fa927898fa937978fff00101fff01101faa23609fba13608fe801209ffd01209ffc0012afd80149afff00101fef01101;
assign testcases[848] = 512'hfab32787fab27787fe702788fe802688fa927898fa937978fff00001fff01101fba23609fba13608fe801209ffd01209ffc0012afd80149afff00101fef00101;
assign testcases[849] = 512'hfef00112fef01112fff00122fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00005fff00015fff00001fff00000;
assign testcases[850] = 512'hfef00122fef01122ffe00223fff00223fef01223fef01223fff00000fff00000fef00104fef00104fff00003fff00103fff00015fff00125fff00001fff00000;
assign testcases[851] = 512'hfdf10233fdf01233ffe01233ffe01233fee02233fee12223fff00000fff00000fef01104fef01204ffe00104fff00104fff00016ffe00135fff00001fff00000;
assign testcases[852] = 512'hfdf11233fdf12233ffe01334ffe01233fee12234fee12334fff00000fff00000fde01205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00001;
assign testcases[853] = 512'hfde11333fde12333ffd01334ffd01334fde12344fde12334fff00000fff00000fde11205fde01205ffd00104fff00104fff00016ffe00136fff00001fff00001;
assign testcases[854] = 512'hfde11344fde13344ffc01444ffd01344fdd13455fdd13445fff00000fff00000fde11305fde11305ffd00105fff01105fff00117fed00247fff00001fef00001;
assign testcases[855] = 512'hfcd21454fcd14454ffc01445ffc01455fdc14455fdd24545fff00000fff00000fdd11306fcd12306ffc00106fff01106ffe00117fec01257fff00001fef00001;
assign testcases[856] = 512'hfcd21465fcd14465ffb01556ffc01455fcc14566fcc25556fff00000fff00000fcd12306fcd12406ffc01106ffe01106ffe00128feb01268fff00001fef00001;
assign testcases[857] = 512'hfcd21565fcd25565fea01566feb01466fcb15676fcb25656fff00000fff00001fcc12407fcc12407ffb01107ffe01207ffe00128feb01368fff00001fef00001;
assign testcases[858] = 512'hfcc21575fbc25575fea02667fea02566fcb15677fcb26767fff00000fff00001fcc12407fcc12507ffb01107ffe01207ffd00129fda01379fff00001fef00001;
assign testcases[859] = 512'hfbc32676fbc26676fe902667fea02577fba26787fba26767fff00000fff00001fbb22507fcc12507ffa01107ffe01208ffd00129fda01379fff00001fef00001;
assign testcases[860] = 512'hfbc32676fbc26686fe902677fea02577fba26787fba37877fff00000fff00001fbb22508fbb12508fea01108ffe01208ffd0012afd901489fff00001fef00001;
assign testcases[861] = 512'hfbb32686fbb27786fe802678fe902677fb926898fb937878fff00000fff00001fbb23508fbb13508fe901208ffe01208ffd0012afd80148afff00001fef00001;
assign testcases[862] = 512'hfef00112fef01112fff00122fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00005fff00025fff00001fff00000;
assign testcases[863] = 512'hfef10123fef01122ffe00223fff00223fef01223fef01223fff00000fff00000fef00104fef00104fff00003fff00103fff00015fff00125fff00001fff00000;
assign testcases[864] = 512'hfdf10233fdf02233ffe01233ffe01233fee02234fee12223fff00000fff00000fef01104fef01204ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[865] = 512'hfdf11233fdf12233ffd01334ffe01233fee12334fee12334fff00000fff00000fde11205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00001;
assign testcases[866] = 512'hfde11333fde12343ffd01334ffe01334fde12344fde12334fff00000fff00000fde11205fde01205ffe00105fff00104fff00016ffe00136fff00001fff00001;
assign testcases[867] = 512'hfde11344fde13344ffc01445ffd01344fdd13455fdd13445fff00000fff00000fdd11306fde11305ffd00105fff01105fff00117fed00257fff00001fef00001;
assign testcases[868] = 512'hfcd21454fcd14454ffc01445ffc01455fdc14455fdd24545fff00000fff00000fdd11306fdd12306ffc00106fff01106ffe00118fec01257fff00001fef00001;
assign testcases[869] = 512'hfcd21565fcd14565ffb01556ffc01455fcc14566fcc25656fff00000fff00000fcc12406fcd12406ffc01106ffe01106ffe00128feb01368fff00001fef00001;
assign testcases[870] = 512'hfcd21565fcd25565ffa01556feb01466fcb15676fcb25656fff00000fff00001fcc12407fcc12407ffb01107ffe01207ffe00128feb01368fff00001fef00001;
assign testcases[871] = 512'hfcc21565fcc25575fea02566feb02566fcb15677fcb26767fff00000fff00001fcc12407fcc12507ffb01107ffe01207ffd00129fda01379fff00001fef00001;
assign testcases[872] = 512'hfbc32676fbc26676fe902667fea02577fba26787fba36767fff00000fff00001fbb22507fbb12507ffa01107ffe01208ffd00129fd901379fff00001fef00001;
assign testcases[873] = 512'hfbc32676fbc26686fe902677fea02577fba26787fba37877fff00000fff00001fbb22508fbb12508fea01108ffe01208ffd0012afd901489fff00001fef00001;
assign testcases[874] = 512'hfbb32686fbb27686fe802678fe902677fb926898fb937878fff00000fff00001fbb23508fbb13508fe901108ffe01208ffd0012afd80148afff00001fef00001;
assign testcases[875] = 512'hfef00112fef01112fff00122fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00005fff00015fff00001fff00000;
assign testcases[876] = 512'hfef10123fef01122ffe00223fff00223fef01223fef01223fff00000fff00000fef00104fef01104fff00004fff00103fff00015fff00125fff00001fff00000;
assign testcases[877] = 512'hfef10233fdf02233ffe01233ffe01233fee02234fee12223fff00000fff00000fef01104fef01204ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[878] = 512'hfdf11233fdf12233ffe01334ffe01233fee12334fee12334fff00000fff00000fde11205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00001;
assign testcases[879] = 512'hfde11333fde12333ffd01334ffe01334fde12334fde12334fff00000fff00000fde11205fde01205ffe00105fff00104fff00016fed00136fff00001fff00001;
assign testcases[880] = 512'hfde11344fde13344ffc01445ffd01344fdd13445fdd13435fff00000fff00000fdd11305fde11305ffd00105fff01105fff00117fed00247fff00001fef00001;
assign testcases[881] = 512'hfcd21444fcd14454ffc01445ffc01455fdc14555fdc24545fff00000fff00000fcd11306fdd11306ffc00106fff01106ffe00117fec01257fff00001fef00001;
assign testcases[882] = 512'hfcd21555fcd14555ffb01556ffc01455fcc14566fcc25646fff00000fff00000fcd12406fcd12406ffc01106ffe01106ffe00118feb01358fff00001fef00001;
assign testcases[883] = 512'hfcd21565fcd25565ffa01556ffb01466fcb15666fcb25656fff00000fff00001fcc12407fcc12407ffb01107ffe01207ffe00128feb01368fff00001fef00001;
assign testcases[884] = 512'hfbc21565fcc25575fea02566feb02566fcb15677fcb26767fff00000fff00001fcc12407fcc12507ffb01107ffe01207ffd00129fda01378fff00001fef00001;
assign testcases[885] = 512'hfbc32676fbc26676fe902667fea02567fba26787fba26767fff00000fff00001fbb22507fbb12507ffa01107ffe01208ffd00129fd901379fff00001fef00001;
assign testcases[886] = 512'hfbb32676fbb26676fe902677fe902677faa26788faa37867fff00000fff00001fab22508ebb13508fea01108ffe01208ffd0012afd901489fff00001fef00001;
assign testcases[887] = 512'hfbb32786fbb27786fe802778fe902677fb926898fb937878fff00000fff00001fba23508fbb13608fe901208ffe01208ffd0112afd80148afff00001fef00001;
assign testcases[888] = 512'hfef00112fef01112fff00112fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00005fff00015fff00001fff00000;
assign testcases[889] = 512'hfef10223fef01223ffe01223fff01223fef01223fef11223fff00000fff00000fef01104fef01104fff00004fff00103fff00016fff00125fff00001fff00000;
assign testcases[890] = 512'hfdf10233fdf12233ffe01233ffe01233fee02234fee12224fff00000fff00000fdf01205fef01204ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[891] = 512'hfde11233fde12233ffd01334ffe01234fee12334fee12334fff00000fff00000fde11205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[892] = 512'hfde11333fde12343ffd01334ffd01334fde12344fde13334fff00000fff00000fde11205fde01205ffd00105fff00104fff00016fed00246fff00001fff00001;
assign testcases[893] = 512'hfde11444fde13444ffc01445ffd01344fdd13455fdd13445fff00000fff00000fdd11306fdd11306ffd00105fff01105fff00117fed00247fff00001fef00001;
assign testcases[894] = 512'hfcd21454fcd14454ffb01455ffc01455fdc14555fdc24545fff00000fff00000fcd12306fcd12306ffc00106fff01106ffe00118fec01257fff00001fef00001;
assign testcases[895] = 512'hfcd21555fcd15565ffb01556ffb01456fcc14566fcc25656fff00000fff00000fcc12407fcc12406ffc01106ffe01106ffe00128feb01368fff00001fef00001;
assign testcases[896] = 512'hfcc21565fcc25565fea02566feb02566fcb15676fcb25656fff00000fff00001fcc12407fcc12407ffb01107ffe01207ffe00129fea01368fff00001fef00001;
assign testcases[897] = 512'hfbc31666fbc26676fe902667fea02567fbb16677fbb26767fff00000fff00001fbb22507fcc12507ffa01107ffe01208ffd00129fda01379fff00001fef00001;
assign testcases[898] = 512'hfbc32676fbc26676fe902667fea02577fba26787fba37767fff00000fff00001fbb22508fbb12508ffa01108ffe01208ffd0012afd901479fff00001fef00001;
assign testcases[899] = 512'hfbb32676fbb27776fe902678fe902677fba26788fba37868fff00000fff00001fbb23508fbb13508fea01108ffe01208ffd0012afd90148afff00001fef00001;
assign testcases[900] = 512'hfbb32786fbb27787fe802778fe902678fa927898fa937878fff00000fff00001fba23608fba13608fe901209ffd01209ffc0112afd80148afff00001fef00001;
assign testcases[901] = 512'hfef00112fef01112fff00122fff00122fef01113fef01113fff00000fff00000fef00104fef00104fff00003fff00003fff00005fff00115fff00001fff00000;
assign testcases[902] = 512'hfef10223fef01223ffe01223fff01223fef01223fef11223fff00000fff00000fef01104fef01104fff00004fff00103fff00016fff00125fff00001fff00000;
assign testcases[903] = 512'hfdf10233fdf12233ffe01233ffe01233fee02234fee12224fff00000fff00000fdf01205fef01205ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[904] = 512'hfde11333fde12233ffd01334ffe01334fee12334fee12334fff00000fff00000fde11205fde01205ffe00104fff00104fff00016ffe00136fff00001fff00000;
assign testcases[905] = 512'hfde11333fde12343ffd01334ffd01334fde13344fde13334fff00000fff00000fde11205fde11205ffd00105fff00105fff00017fed00236fff00001fff00001;
assign testcases[906] = 512'hfde11444fde13444ffc01445ffd01345fdd13455fdd14445fff00000fff00000fdd11306fdd11306ffd00105fff01105ffe00117fed01247fff00001fef00001;
assign testcases[907] = 512'hfcd21454fcd14454ffb01555ffc01455fdc14555fcc24546fff00000fff00000fcd12306fcd12406ffc01106fff01106ffe00118fec01257fff00001fef00001;
assign testcases[908] = 512'hfcd21555fcd25565ffb01556ffb01456fcc15566fcc25656fff00000fff00000fcc12407fcc12407ffb01106ffe01107ffe00128feb01368fff00001fef00001;
assign testcases[909] = 512'hfcc21565fcc25565fea02566feb02566fcb15676fcb26757fff00000fff00001fcc12407fcc12407ffb01107ffe01207ffe00129fea01368fff00001fef00001;
assign testcases[910] = 512'hfbc32666fbc26676fe902667fea02567fbb26777fbb26767fff00000fff00001fbb22507fcc12507ffa01107ffe01208ffd00129fda01379fff00001fef00001;
assign testcases[911] = 512'hfbc32676fbc26676fe902667fea02577fba26787fba37867fff00000fff00001fbb22508fbb13508ffa01108ffe01208ffd0012afd901479fff00001fef00001;
assign testcases[912] = 512'hfbb32776fbb27786fe802778fe902677fba26788fba37878fff00000fff00001fbb23508fbb13608fea01208ffe01208ffd0012afd90148afff00001fef00001;
assign testcases[913] = 512'hfbb32786fbb27787fe802778fe902678fb927898fa937878fff00000fff00001fba23608fba13608fe901208ffe01209ffd0112afd80148afff00001fef00001;
assign testcases[914] = 512'hfef00123fef01123ffd01334ffd01334fef01123fef01123fdd12313fed12313fef00104fef00104ffe00105fff00104fff00016fff00125fed01303fde12203;
assign testcases[915] = 512'hfdf00123fef01123ffd01334ffd01334fef01123fef01123fdd12313fed12313fef00104fef00104ffe00105fff00105fff00016fff00125fed01303fde12203;
assign testcases[916] = 512'hfdf00223fdf01123ffd01334ffd01334fef01123fef01123fdd12313fed12313fef00105fef00104ffe00105fff00105fff00016fff00125fed01303fde12203;
assign testcases[917] = 512'hfdf00223fdf01123ffd01334ffd01334fef01123fef01223fdd12313fed12313fef00105fef00104ffe00105fff00105fff00016fff00125fed01303fde12203;
assign testcases[918] = 512'hfef10113fef01112ffd01324ffd01324fef11113fef01112edd53313fdc65414fef00104fef00104ffe00104fff00104fff00005fff00015fed02304fde13303;
assign testcases[919] = 512'hfef00123fef01123ffd01334ffd01334fef01123fef01113fdd23314fdc24415fef00104fef00104ffe00104fff00104fff00005fff00025fed02404fde13303;
assign testcases[920] = 512'hfef00123fef01123ffd01334ffd01334fef01123fef01113fdd23314fdc24415fef00104fef00104ffe00104fff00104fff00005fff00025fed02404fde13303;
assign testcases[921] = 512'hfef10123fef11123ffd01334ffe01334fef11123fef01113fdd43314fdc54415fef10104fef00104ffe00104fff00104fff00005fff00025fed13404fde23303;
assign testcases[922] = 512'hfef00123fef01123ffd01334ffd01334fef01123fef01113edd23314fdc24515fef00104fef00104ffe00104fff00104fff00005fff00025fed02404fde13303;
assign testcases[923] = 512'hfbc32636fcc26636fe902748fea02647fba26737fbb26837fff00000fff00000fbb23608fbb23608ffa01208ffe01208ffd0111afd901439fff00001fef00001;
assign testcases[924] = 512'hfbc32736fcc26636fe903748fea02647fba27737fba37837fff00000fff00000fbb23608fbb23608ffa01208ffe01208ffd0111afd90143afff00001fef00001;
assign testcases[925] = 512'hfcd215b4fcd144b4fe814a69fe913858fdd155c5fdc255c5fff00000fff00000fcd12406fcd12406fe901209ffe01209ffe00138fec013c8fff00001fef00001;
assign testcases[926] = 512'hfcd21434fcd14434fe714949fe913848fdd15535fdc24535fff00000fff00000fcd12406fcd12406fe901209ffe01209ffe00118fec01337fff00001fef00001;
assign testcases[927] = 512'hfcd31555fcd25554fe814a69fe913858fcc25555fcc25646fff00000fff00000fcc22407fcc13507fea01209ffe02309ffe00118feb01358fff00001fef00001;
assign testcases[928] = 512'hfcd21535fcd25434fe713959fe913858fcc15545fcc25536fff00000fff00000fcc12407fcc12407fe901209ffe01209ffe00118feb01338fff00001fef00001;
assign testcases[929] = 512'hfcd215f4fdd144f4fe814a69fe913868fdd155f5fdd255f5fff00000fff00000fcd12406fcd12406fea01209ffe01209ffe00148fec013f8fff00001fef00001;
assign testcases[930] = 512'hfcd21434fcd14434fe713949fe913848fdd14535fdc24535fff00000fff00000fcd12406fcd12406fe901208ffe01209ffe00118fec01337fff00001fef00001;
assign testcases[931] = 512'hfcd32665fcd26565fe814959fe913858fcc26666fcc26656fff00000fff00000fcc22407fcc23507fea01208ffe01209ffe00129feb01368fff00001fef00001;
assign testcases[932] = 512'hd9a53a67daa39967fd215f7dfd414c7ce9839a79d984ab69fff00000fff00001d993480ad992590afe51230cffc0240cffc0122cdb60267bfff00101fef00001;
assign testcases[933] = 512'hfaa42847fbb38737fd314c5cfe514a5cfa828948fa839a39fff00000fff00000fa92470afa924709fe60130bffd0230cffc0111bfc60154bfff00001fef00001;
assign testcases[934] = 512'hfaa42867fbb27767fd414dadfe514bbcfa928869fa938959fff10010fff10010fa92370afa92470afe61130cffd1230cffc0112bfd70156bfff00001fef00001;
assign testcases[935] = 512'hfcd31535fcd25535fe813848fea13748fcc15646fcc25636fff00000fff00000fcc22407fcc13507ffa01208ffe01208ffe00118feb01348fff00001fef00001;
assign testcases[936] = 512'hfcd31545fcd25545fe813858fea13758fcc15646fcc25646fff00000fff00000fcc22507fcc13507ffa01208ffe01208ffe00119feb01348fff00001fff00001;
assign testcases[937] = 512'hfcd32655fcd26555fe814958fea13858fcc26666fcc26756fff00000fff00000fcc23507fcc23507ffa01208ffe01208ffe00119feb01358fff00001fef00001;
assign testcases[938] = 512'hfcd21564fcd24464fe913747fea12647fdd15565fdc25575fff00000fff00000fcd12406fcd12406ffb01207ffe01207ffe00128fec01378fff00001fff00000;
assign testcases[939] = 512'hfcd32655fcd26555fe913958fea13758fcc26656fcc37746fff00000fff00000fcc23507fcc23507ffa01208ffe01208ffe01119feb01458fff00001fef00001;
assign testcases[940] = 512'hfcd32655fcd26555fe913858fea13757fcc26666fcc36756fff00000fff00000fcc23507fcc23507ffb01208ffe01208ffe00119feb01358fff00001fef00001;
assign testcases[941] = 512'hfcd32655fcd26555fe913958fea13758fcc26656fcb37746fff00000fff00000fcc23507fcc23507ffa01208ffe01208ffe01119fea01459fff00001fff00001;
assign testcases[942] = 512'hfcd32645fcd26545fe913848fea13747fcc26656fcb36746fff00000fff00000fcc23507fcc13507ffa01208ffe01208ffe00119fea01459fff00001fff00001;
assign testcases[943] = 512'hfbb42886fbc38786fe413bacfe513aacfcb27876fcc38966ecc24455fdb24455fbb23708fbb24708fe70120cffd0130cffe01128feb01468fdc02405ecc13314;
assign testcases[944] = 512'hfbb21667fbb14566fe413a9cfe513a9cfcb14566fcb14456ecb35555fdb25555fbb12408fbb12408fe70120cffd0130bffe00118feb01268fdb13505ecc15404;
assign testcases[945] = 512'hfbc21655fcc14555fe613a7afe71397afcc14545fdd13445edd36533fdc36533fcc12407fcc12407fe901209ffe01309ffe00117fec01247fed13503edd15503;
assign testcases[946] = 512'hfcc31555fcd25455fe714a6afe814a6afdc14455fdd24445edd24443fdd24443fcc12407fcc12407fe90120affe0130affe00118fec01247fec03404fdd14413;
assign testcases[947] = 512'hfcc32656fcc25555fe614b6bfe714a6bfcc15556fcc25546edd24453fdc24443fcc22408fcc12508fe80120affe0230affe00118fec01248fec03404edd14413;
assign testcases[948] = 512'hfcc315b6fcd245a5fe714a8afe82498afdc244a6fdd24476edd24373fdd24463fcd22307fcd12407fe91120affe1220afff00127fed01287fed02414edd14313;
assign testcases[949] = 512'hfcd31555fcd25545fe914969fe914969fdd14445fdd24435ede23353fed13353fcc22407fcc12407ffa11209ffe12209ffe00118fec01247fed02303fde13313;
assign testcases[950] = 512'hfcd31535fcd24545fe813959fe914959fdd15435fdd24435ede33343fed33343fcc12407fcc12407ffa11209ffe12209ffe00118fec01237fed02303fde23313;
assign testcases[951] = 512'hfde31424fde24334ffa13747ffb13747fde13324fde23324fee12232fee12232fdd12306fdd12306ffc11207fff11207fff00017ffe00226fee01202fee02202;
assign testcases[952] = 512'hfde21434fde13334ffb13747ffb13747fee13334fee13324fee12232fee12232fde11205fde11305ffc01107fff01206fff00016ffe00126ffe01202fee02202;
assign testcases[953] = 512'hfab32767fbb25667fe414b7cfe514b7cfcb15667fcb25657ecc35544edc25544fbb12508fbb12508fe70120bffd0130bffe00119feb01248edb13505ecc15504;
assign testcases[954] = 512'hfcc32645fcd26545fe913848fea13747fcc26646fcb36747fff00000fff00000fcc23507fcc13507ffa01208ffe01208ffe00119fea01449fff00001fff00001;
assign testcases[955] = 512'hfcc42655fcd27655fe913858fea13757fcc27666fcb37756fff00000fff00000fcc23507fcc23607ffa01208ffe01208ffe01119fea01459fff00001fff00001;
assign testcases[956] = 512'hfde31534fde25434ffb13746ffc13636fdd15545fdd25635fff00000fff00000fdd22406fdd12406ffc01106fff01206ffe00118fec01347fff00001fff00000;
assign testcases[957] = 512'hfbb42867fbc38766fe713a6afe813869fba28878fba49968fff00000fff00000fba34609fba24709fe901209ffe01209ffd0112afd90157afff00001fef00001;
assign testcases[958] = 512'hfab42868fbb27767fe515c8cfe615c8cfba26767fba36748ecc34474fdc25474fba23609fba23609fe71230cffd1230cffd00119fda01359fdc13504ecc15414;
assign testcases[959] = 512'hfde11314fde12313fe502a5bfe80285afdd13515fde13414fff00001fff00001fde11406fde11406fe90120affe01209ffe00108fed01317fff00101fef01101;
assign testcases[960] = 512'hfde11314fde12313fe502a5cfe80285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[961] = 512'hfde11314fde12313fe502a5cfe80285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[962] = 512'hfde11314fde12313fe502a5cfe80285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[963] = 512'hfde11314fde12313fe502a6cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[964] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[965] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[966] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[967] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[968] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[969] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[970] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00109fed01328fff00101fef01101;
assign testcases[971] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[972] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00109fed01328fff00101fef01101;
assign testcases[973] = 512'hfde11314fde12313fe502a6cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00109fed01328fff00101fef01101;
assign testcases[974] = 512'hfde11314fde12313fe502a6cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00109fed01328fff00101fef01101;
assign testcases[975] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00109fed01328fff00101fef01101;
assign testcases[976] = 512'hfde11314fde12313fe502a6cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00109fed01328fff00101fef01101;
assign testcases[977] = 512'hfde11314fde12313fe502a6cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00109fed01328fff00101fef01101;
assign testcases[978] = 512'hfde11314fde12313fe502a5cfe70285afdd13515fde13414fff00001fff00001fdd11406fde11406fe90120affe01209ffe00108fed01328fff00101fef01101;
assign testcases[979] = 512'hfde11313fdf12313fe70294afe902749fde13415fee12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01328fff00101fef00001;
assign testcases[980] = 512'hfde11313fde12313fe70294afe902849fde13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01328fff00101fef00001;
assign testcases[981] = 512'hfde11313fde12313fe70294bfe902849fde13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[982] = 512'hfde11313fde12313fe70294afe902849fdd13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[983] = 512'hfde11313fdf12313fe70294bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[984] = 512'hfde11313fde12313fe70294bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[985] = 512'hfde11313fde12313fe70295bfe902849fde13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[986] = 512'hfde11313fde12313fe70294bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[987] = 512'hfde11313fde12313fe70295bfe902849fdd13415fde12314fff00001fff00001fde11306fde11406fea01209ffe01208fff00108fed01328fff00101fef00001;
assign testcases[988] = 512'hfde11313fde12313fe60295bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[989] = 512'hfde11313fde12313fe70295bfe902849fdd13415fee12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[990] = 512'hfde11313fde12313fe60295bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306fea01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[991] = 512'hfde11313fde12313fe60295bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306fea01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[992] = 512'hfde11313fde12313fe60295bfe802849fdd13415fde12314fff00001fff00001fde11306fde11306fea01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[993] = 512'hfde11313fde12313fe70294bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01217fff00101fef00001;
assign testcases[994] = 512'hfde11313fde12313fe70295bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01227fff00101fef00001;
assign testcases[995] = 512'hfde11313fde12313fe60295bfe902849fdd13415fee12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[996] = 512'hfde11313fde12313fe60295bfe802849fdd13415fde12314fff00001fff00001fde11306fde11306ffa01209ffe01208fff00108fed01228fff00101fef00001;
assign testcases[997] = 512'hfde11313fde12313fe70295bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306fea01209ffe01208fff00108fed01227fff00101fef00001;
assign testcases[998] = 512'hfde11313fde12313fe60295bfe902849fdd13415fde12314fff00001fff00001fde11306fde11306fea01209ffe01208fff00108fed01227fff00101fef00001;
assign testcases[999] = 512'hfdf10213fdf01213fe901749fea01638fee12315fee12314fff00000fff00000fde11306fde01306ffb00108fff01207fff00108ffe00217fff00101fef00001;



gasId_tnn1_tnnpar dut (.features(features),.prediction(prediction));

integer i,j;
initial begin
    features = testcases[0];
    for(i=0;i<TEST_CNT;i=i+1) begin
        features = testcases[i];
        #period
        /* $display("%h",features); */
        /* $display("%b",dut.hidden); */
        for(j=0;j<CLASS_CNT;j=j+1) begin
            $write("%d ,",dut.scores[j]);
        end
        $display("");
        $display("%d",prediction);
    end
end

endmodule
