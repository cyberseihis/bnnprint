
















module Har_bnn1_bnnpaarx #(

parameter FEAT_CNT = 12,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 4448'h0064008700560086004f00790068007800520077005900760049007500490074004a007200630071005c00700044006f0045006e0061006d0042006c0045006b003c006a0055006900570067005a0066003b00650046006200420060004e005f003c005e0054005d0046005b003b00580036005400220053001d0053003f0052003e0051002b0051004b0050002b00500047004f004d004e0040004d004a004c0043004c001e004b003b00480024004800330047002a004400340043003c00420032004100330040002e00400031003d001c003a00340039002e003800210038002900370027003700280036002c003500260035001d0035002900300026002f0027002d0020002d0023002c0019002b0028002a0024002a001b00280023002500200025001c002500210022001b002200180020001e001f001f0041002a003f001a003e0018003d0032003a0030003900360038002e003700280035001d00310024002f002d002e0021002d0029002b001a002b0026002a002500280020002400310034002200330018003200270030001d002f00230029001c0027001b00250019002400180019001c002c001b002600030015001e0023001a002200110014001c001e00040016000e0012000a0010000500080002000600000001001d0020001a001b0009000f0007000b00180021001300170001000c000c000d0019001f00070017000800110004000a0006000e00030009000b00130002001200100016000f0015000500140000000d ;
localparam YMAP = 640'h00a1007c008800970081008e0095008a00930083009800850084008b009f008f0080008c007b009c009100940090009b007f0089007d0073009a009e008d007a009d007e00a2009200960099008200a0;
localparam ADDCNT = $bits(PAAR0) / 32;
localparam FULLCNT = ADDCNT + (FEAT_CNT * 2);
localparam PAAR1 = 3296'h00a800b000a900af00a700ae00aa00ad00a600ac00a000ab00a100a5009d00a4009a00a3009e00a20099009f008c009c008e009b0093009800950097008d009600900094008f0092008a00910081008b0086008900850088008400870084008600830085008200830075008200600081007e007f007c007f0065007e0078007c0076007900670071005d006f00620063005f0061003b005e0023005800390057003c0056004b0054003d004a0019004900040037001100290001001900130018007a00800075007d0079007b000c0078006f00760013007100420067000000650017004d002e004c0014003b0007003a000a00360074007700690073006d0072006a0070006c006e0068006b00640066005f00630003006200480061002b0060005d005e0047004f00330045004300440002003c002700300008002d0020002a001c001f000b001d0005001b005a005c0058005b0032005900410057003400560028004b0025003f002900390012002f00060024000e001a0040005500210054000f002c0015002200520053005000510035003e001e002600090010 ;
localparam YMAP1 = 96'h00b300b500b600b400b200b1;
localparam ADDCNT1 = $bits(PAAR1) / 32;
localparam FULLCNT1 = ADDCNT1 + (HIDDEN_CNT * 2);
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[FEAT_CNT+i] = -feature_array[i];
endgenerate

integer j;
generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam op1 = PAAR0[i*32+:16];
    localparam op2 = PAAR0[i*32+16+:16];
    localparam nodeloc = (2 * FEAT_CNT) + i;
    assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    assign hidden[i] = node[YMAP[i*16+:16]] >= 0;
end
endgenerate

/* initial begin */
/*     #10 */
/*     for(j=0;j<FULLCNT;j=j+1) */
/*         $display("%d | %d", j, node[j]); */
/* end */

wire unsigned [SUM_BITS-1:0] xnode [FULLCNT1-1:0];

generate
    for(i=0;i<HIDDEN_CNT;i=i+1)
        assign xnode[i] = hidden[i];
    for(i=0;i<HIDDEN_CNT;i=i+1)
        assign xnode[HIDDEN_CNT+i] = hidden_n[i];
for(i=0;i<ADDCNT1;i=i+1) begin
    localparam op1 = PAAR1[i*32+:16];
    localparam op2 = PAAR1[i*32+16+:16];
    localparam nodeloc = (2 * HIDDEN_CNT) + i;
    assign xnode[nodeloc] = xnode[op1] + xnode[op2];
end
for(i=0;i<CLASS_CNT;i=i+1) begin
    assign scores[i*SUM_BITS+:SUM_BITS] = xnode[YMAP1[i*16+:16]];
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
