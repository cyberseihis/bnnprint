module binaccum #(
    parameter N = 4 // Number of elements to add
)(
    input clk,             // Clock input
    input rst,             // Reset input
    input put,
    input unsigned data_in,  // Input data
    output reg unsigned [$clog2(N+1)-1:0] acc
);

always @(posedge clk or posedge rst) begin
    if (rst) begin
        acc <= 0;
        $display(N);
    end else if (!put) begin
        acc <= acc+data_in;
        $display("tt %t",$time);
        /* $display("ba %d",acc); */
    end
end

endmodule
