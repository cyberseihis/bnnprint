`timescale 1us/1ns









module tbgasId_bnn1_bnnseq #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)();

  
  reg [FEAT_BITS*FEAT_CNT-1:0] sample;
  wire [FEAT_BITS*FEAT_CNT-1:0] testcases [TEST_CNT-1:0];
  reg rst;
  reg clk;
  parameter Nsperiod=50000;
  localparam period=Nsperiod/500;
  localparam halfPeriod=period/2;


assign testcases[0] = 512'h10000fef10000fff41000fff50000fff20000fff30000fff30000fef30000fef10000fff10000fff21000fff21000fff21000fff21100fff21000fef21000fef;
assign testcases[1] = 512'h10100fef10100fff41000fff50000fff20000fff30000fff30000fef40000fef10100fff10110fff21100fef21000fef22100fff22100fff21000fef21000fef;
assign testcases[2] = 512'h10110fef20100fff51000fff50000fff30000fff40000eff40100fef40100fef10110fff10111fef31110fef32100fef32100eff32100eff22100fef22100fef;
assign testcases[3] = 512'h10111fef20110fff51100fff50000fff30000fff40000eff40100fef40100fef10111fff10111fef31110fef32110fef32200eff32200eff22110fef22100fef;
assign testcases[4] = 512'h20110fef20110eff52100fff51000fff30000fff40000eff40100fef40100fef20111eef20111eef32110fef32110fef33200eff43200dff22110fef32100fef;
assign testcases[5] = 512'h20220edf30210eef52100eff61000fff40100fff50100dff50100edf50100edf21221eef21221edf32210eef33110eef44210dff44310cff33110fdf33101fdf;
assign testcases[6] = 512'h30221edf30210def63100eff61000fff50100fff60100cff50210edf50110edf31221def31232ddf42211eef43210eef54310cff54310bff33210edf33201edf;
assign testcases[7] = 512'h30231ddf30320def63100def61000fff50100fff60100bff50210edf50210edf31331ddf31332ddf43211edf44210edf55310cff55410bef44210edf44201edf;
assign testcases[8] = 512'h30331ddf40320def64100def71000fff60100fff70100bff60210ddf60210ddf31332ddf31332cde43221ddf44220ddf66310bef66410aef45221edf45201dcf;
assign testcases[9] = 512'h30331ddf40320cef74100cef71000fff60100eff70100aef60210dcf60211dcf41332cdf41342cce53321ddf55220ddf66310aef764109ef45221dcf45301dcf;
assign testcases[10] = 512'h40341dce40420cef74100cef71000eff70100eff801009ef60210ccf60211ccf41342cdf41442cce54321ccf55321ccf774109ef774108ef56321dcf56311dcf;
assign testcases[11] = 512'h40341ccf50430cef75100bef81000eff70100eff801008ef70211ccf70211ccf41442cdf41443cce64321ccf55321ccf774109ef875107ef56321ccf56311cbf;
assign testcases[12] = 512'h40451cce50430cef85200bef81000eff70100eff901008ef70311bbf70211bcf41442bde51453bce64321bcf66321bcf884108ef885106ef56321cbf56311cbf;
assign testcases[13] = 512'h40451cce50430bdf85200adf81000eff80100eff901007ef70311bbf70311bbf51452bdf51453bce65321bbf66321bcf884107ef885106ef67321bbf57311bbf;
assign testcases[14] = 512'h10000fef10000fff41000fff50000fff20000fff30000fff30000fef30000fef10000fff10000fff21000fff21000fff21100fff21100fff21000fef21000fef;
assign testcases[15] = 512'h10110fef10100fff51000fff50000fff30000fff30000fff40100fef40000fef10110fff10110fef31100fef31100fef32100fff32100eff21100fef21100fef;
assign testcases[16] = 512'h10110fef20110fff51000fff50000fff30000fff40000eff40100fef40100fef10110fff10111fef31110fef32110fef32100eff32200eff22110fef22100fef;
assign testcases[17] = 512'h20110fef20110eff52100fff50000fff40000fff40000eff40100fef40100fef20111fff20111eef31110fef32110fef33200eff43210dff32110fef32100fef;
assign testcases[18] = 512'h20110fef20210eff52100eff60000fff40100fff50100dff40100fef40100fef20221eef21221eef31210fef32110fef43210dff43310dff32110fef32100fdf;
assign testcases[19] = 512'h20220edf30210eef62100eff61000fff50100fff50100cff50210edf50110edf21221eef21221edf42211eef43210eef44310cff54310cff33210edf33201edf;
assign testcases[20] = 512'h30221edf30320def63100def61000fff50100fff60100bff50210ddf50210edf31231def31332dde42221edf43210edf54310cff64410bef43220edf43201edf;
assign testcases[21] = 512'h30331ddf30320def73100def71000fff60100fff70100bff60210dcf60211ddf31331def31332ddf53321ddf43220ddf65410bef65410aef44221ddf44311dcf;
assign testcases[22] = 512'h30331ddf40320def73100cef71000eff60100eff70100aef60210dcf60211dcf31331ddf31332cde53321ddf54321ddf66410aef764109ef44321dcf44311dcf;
assign testcases[23] = 512'h30331ddf40320cef74100cef71000eff70100eff801009ef60311ccf70211ccf41342cdf41342cce53321ccf54321ccf76410aef765108ef55321dcf55311dcf;
assign testcases[24] = 512'h40341dcf40420cef84200bef81000eff70100eff801009ef70311cbf70311ccf41442cdf41442cce64421ccf55321ccf774109ef865107ef55321ccf55311cbf;
assign testcases[25] = 512'h40341dcf40420cef85200aef81000eff80100eff901107ef70311bbf70311bbf41442cdf41443cce64421bcf65321bcf875108ef875206ef56321cbf56411cbf;
assign testcases[26] = 512'h40441ccf50430cef85200adf81100eff80110dff901107ef70311bbf70311bbf41442cdf51453bce64431bbf66431bbf875107ef976206ef66421bbf66411bbf;
assign testcases[27] = 512'h40451cce50430bdf95200adf91100dff80110dffa01106ef80311aaf80311abf51442bdf51453bce75431abf66431abf885107ef986205df67421baf67411baf;
assign testcases[28] = 512'h10000fef10000fff41000fff50000fff20000fff30000fff30000fef30000fef10000fff10000fff21000fff21000fff21000fff21100fff21000fef21000fef;
assign testcases[29] = 512'h10110fef10100fff51000fff50000fff30000fff30000fff40000fef40000fef10110fff10110fef21100fef21100fef22100fff32100eff21000fef21100fef;
assign testcases[30] = 512'h10110fef20110fff51000fff50000fff30000fff40000eff40100fef40100fef10110fff10111fef31110fef31110fef32100eff32200eff22110fef22100fef;
assign testcases[31] = 512'h20110fef20110eff52100fff50000fff30000fff40000eff40100fef40100fef20111fff20111eef31110fef32110fef33200eff43200dff22110fef22100fef;
assign testcases[32] = 512'h20110fef20210eff52100fff61000fff40100fff40100dff40100fef40100fef20221eef20221eef32110fef32110fef43210dff43310dff32110fef32100fdf;
assign testcases[33] = 512'h20220edf30210eef63100eff61000fff40100fff50100cff50100edf50100edf21221eef21221edf42210eef43210eef44310dff54310cff33210edf33201edf;
assign testcases[34] = 512'h30221edf30320def63100eff61000fff50100fff60100cff50210edf50210edf31231def31332ddf42211edf43210edf55310cff55410bff34210edf34201edf;
assign testcases[35] = 512'h30231ddf30320def64100def71000fff50100fff60100bff60210ddf60210ddf31331def31332ddf43221ddf44210ddf55310bff65410aef45210edf45201edf;
assign testcases[36] = 512'h30341ddf40320def74100def71000fff60100eff70100aff60210dcf60211dcf31342ddf31342cde53322ddf54321ddf66410bef66510aef45321dcf45311dcf;
assign testcases[37] = 512'h30331ddf40320cef74100cef71000eff60100eff801009ef60210ccf60211ccf41342cdf41342cce53321ccf55321cdf66410aef764109ef55321dcf55311dcf;
assign testcases[38] = 512'h40341dcf40420cef74200bef81000eff70100eff801009ef70311ccf70211ccf41442cdf41442cce64321ccf55321ccf774109ef775108ef56321ccf56311cbf;
assign testcases[39] = 512'h40341cce50430cdf85200bef81000eff70100eff801008ef70311bbf70211ccf41442cde41443bbe64321ccf66321ccf774109ef875107ef56321cbf56311cbf;
assign testcases[40] = 512'h40441cce50430cef85200adf81000eff80100eff901007ef70311bbf70311bbf41442cdf51453bce65421bcf66321bcf884108ef885106ef57321bbf57411cbf;
assign testcases[41] = 512'h40451cce50430bdf85200adf81100eff80100eff901107ef80311bbf70311bbf51452bdf51453bce65431bbf66421bcf885107ef986206ef67421baf67411baf;
assign testcases[42] = 512'h10000fef10000fff41000fff50000fff20000fff30000fff30000fef30000fef10000fff10000fff21000fff21000fff21000fff21100fff21000fef21000fef;
assign testcases[43] = 512'h10110fef10100fff51000fff50000fff30000fff30000fff40000fef40000fef10110fff10110fef21100fef21000fef22100fff32100fff21000fef21100fef;
assign testcases[44] = 512'h10110fef20110fff51000fff50000fff30000fff40000eff40100fef40100fef10110fff10111fef31110fef32110fef32100eff32200eff22110fef22100fef;
assign testcases[45] = 512'h10110fef20110fff51100fff50000fff30000fff40000eff40100fef40100fef10111fff10111fef31110fef32110fef33200eff33200eff22110fef22100fef;
assign testcases[46] = 512'h20110fef20110eff52100fff50000fff40000fff50100dff40100fef40100fef20111eef21221eef31110fef32110fef33200eff43210dff22110fef32100fef;
assign testcases[47] = 512'h20220edf30210eef62100eff61000fff40100fff50100dff50210edf50110edf21221eef21221ddf32211eef33210eef44310dff44310cff33110fdf33201fdf;
assign testcases[48] = 512'h30231edf30320def63100eff61000fff50100fff60100cff50210edf50210edf31331def31332ddf42211eef43210eef55310cff55410bff33210edf33201edf;
assign testcases[49] = 512'h30331edf30320def63100def71000fff50100fff60100bff60210ddf60210ddf31331def31332ddf43221edf43210edf55310cff65410bef44221edf44201edf;
assign testcases[50] = 512'h30331ddf40320def73100def71000fff60100eff70100aff60210dcf60211dcf41342cdf41442cce43221ddf44220ddf66310bef66410aef44221ecf44211dcf;
assign testcases[51] = 512'h30331ddf40320cef74100cef71000eff60100eff70100aef60210ccf60211ccf41442cdf41442cce53321ddf54221ddf66410aef764109ef45221dcf45311dcf;
assign testcases[52] = 512'h40331ddf40420cef74200bef81000eff70100eff801009ef70311ccf70211ccf41442cdf41442cce54321ccf55321ccf774109ef765108ef55321dcf55311dcf;
assign testcases[53] = 512'h40341dcf40420cef85200bef81000eff70100eff901008ef70311bbf70311bbf41442cdf51443bce54321ccf55321ccf774109ef875108ef56321ccf56311cbf;
assign testcases[54] = 512'h40441cce50430cef85200aef81000eff80100eff901007ef70311bbf70311bbf51452bdf51453bce64321ccf56321ccf784108ef875107ef56321cbf56311cbf;
assign testcases[55] = 512'h40441cce50430cef95200adf91000dff80100dffa01107ef80311abf80311abf51452bdf51553bce64321bbf66321bcf884107ef885106ef57321bbf56311bbf;
assign testcases[56] = 512'h10000fef10000fff41000fff50000fff20000fff30000fff30000fef30000fef10000fff10000fff21000fff21000fff21000fff22000fff21000fef21000fef;
assign testcases[57] = 512'h10110fef10100fff51000fff50000fff30000fff30000fff40100fef40000fef10110fff10110fef21100fef21100fef22100fff32100eff21100fef22100fef;
assign testcases[58] = 512'h10110fef20110fff52000fff50000fff30000fff40000eff40100fef40100fef10110fff10111fef31110fef32110fef33100eff33200eff22110fef22100fef;
assign testcases[59] = 512'h20110fef20110eff52100fff61000fff40000fff40000eff40100fef40100fef20111eef21111eef32110fef32110fef33200eff43200dff32110fef32100fef;
assign testcases[60] = 512'h20110fef20210eff52100eff61000fff40100fff50100dff50100edf50100fef21221eef21221eef32110fef32110fef43210dff43310dff32110fdf32101fdf;
assign testcases[61] = 512'h20220edf30210eef63100eff61000fff50100fff50100cff50210edf50110edf21221eef31221ddf42211eef43210eef44310dff54310cff33210edf33201edf;
assign testcases[62] = 512'h30221edf30320def63100def61000fff50100fff60100cff50210edf50210edf31331def31332ddf42221edf43210eef55310cff55410bff34210edf33201edf;
assign testcases[63] = 512'h30331ddf30320def63100def71000fff60100fff70100bff60210ddf60211ddf31332def31342ddf43221edf44220edf55410bff65410aef44221edf44211edf;
assign testcases[64] = 512'h30331ddf40320def74100cef71000fff60100eff70100aff60210dcf60211dcf41342cdf41442cce53321ddf44220ddf66410bef66410aef45221dcf45311dcf;
assign testcases[65] = 512'h40331ddf40320cef74100cef71000eff60100eff80100aef60310ccf60211ccf41442cdf41442cce54321ddf55321ddf66410aef764109ef45321dcf45311dcf;
assign testcases[66] = 512'h40341ddf40420cef74200bef81000eff70100eff801009ef70311ccf70211ccf41442cdf41442cce54321ccf55321ccf774109ef775108ef56321dcf55311dcf;
assign testcases[67] = 512'h40341dcf40420cef85200bef81000eff70100eff801008ef70311bbf70311bbf41442cdf51453bce54321ccf55321ccf774109ef875108ef56321ccf56311cbf;
assign testcases[68] = 512'h40441cce50430cef85200aef81000eff80100eff901008ef70311bbf70311bbf51452bde51453bce64321ccf66321ccf884108ef885107ef57321cbf56311cbf;
assign testcases[69] = 512'h40441cce50430cef85200adf91000eff80100eff901107ef80311abf80311abf51452bdf51553bce65321bcf66321bcf884108ef885106ef57321bbf57411bbf;
assign testcases[70] = 512'h10000fef10000fff41000fff50000fff20000fff30000fff30000fef30000fef10000fff10000fff21000fff21000fff21000fff21100fff21000fef21000fef;
assign testcases[71] = 512'h10110fef10100fff51000fff50000fff30000fff30000fff40100fef40000fef10110fff10110fef21100fef21100fef32100fff32100eff21100fef21100fef;
assign testcases[72] = 512'h10110fef20110fff51000fff50000fff30000fff40000eff40100fef40100fef10110fff10111fef31110fef31110fef32100eff32200eff21110fef21100fef;
assign testcases[73] = 512'h20110fef20110fff52100fff50000fff40000fff40100eff40100fef40100fef20111eef20111eef31110fef32110fef33200eff43210dff22110fef32100fef;
assign testcases[74] = 512'h20231fef20221eff52100eff60000fff40100fff50100dff50211fdf50111fef21243eef21244eef31221fef32211fef43210dff43310dff32111fdf32200fdf;
assign testcases[75] = 512'h20220edf30210eef62100eff61000fff50100fff60100cff50210edf50110edf21221eef31221ddf42211eef42210eef44310dff54310cff32210edf32201edf;
assign testcases[76] = 512'h30221edf30320def62100def71000fff50100fff60100bff60210ddf60210ddf31331def31332dde42221edf43220edf54310cff54410bff43221edf43201edf;
assign testcases[77] = 512'h30331edf30320def73100def71000fff60100fff70100bff60210dcf60211dcf31331def31332ddf42321ddf43220ddf65410bef65410aef43221edf43311ecf;
assign testcases[78] = 512'h30331ddf40320def73100cef71000eff60100eff80100aef60310ccf60211ccf41332cdf41442cce53321ddf54321ddf66410aef755109ef44321dcf44311dcf;
assign testcases[79] = 512'h30331ddf40320def84200bef81000eff70100eff801009ef70311ccf70311ccf41442cdf41442cce53321ccf54321cdf76410aef765109ef55321dcf55311dcf;
assign testcases[80] = 512'h40341ddf40420cef84200bef81000eff70100eff801008ef70311bbf70311bbf41442cdf41442cce54321ccf55321ccf774109ef765108ef55321cbf55311cbf;
assign testcases[81] = 512'h40341ddf40420cef85200aef81000eff80100eff901108ef80311bbf70311bbf41442cdf51443bce64321ccf55321ccf774108ef875207ef56321cbf56411cbf;
assign testcases[82] = 512'h40441dcf50430cef95200adf91100dff80100eff901107ef80311abf80311abf51442bdf51453bce64421bcf66321bcf885108ef875206ef56421bbf56411cbf;
assign testcases[83] = 512'h40441ccf50430cef96200adf92100dff80100effa01107ef80411abf80311abf51452bdf51553bce65421bbf66321bcf885108ef986206ef67421bbf67411bbf;
assign testcases[84] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff30000fef40000fef00000fff00000fff21000fef21000fff21000fff21000fff21000fef21000fef;
assign testcases[85] = 512'h10000fef10000fff63100eef61000fff30000fff40000dff50100edf50100edf00000fff00000fff42210edf33210eef33200eff33200dff33210edf33200edf;
assign testcases[86] = 512'h00000fff00000fff40200fff40100fff10100fff20100fff30310fef30311fef00000fff00000fff20431fff20321fff10310fff10410fff10321fef10311fef;
assign testcases[87] = 512'h10000fef10000fff74200cef71000eff40100fff50100cff60310ddf60211ddf10000fff00000fff53321ddf44321ddf44310dff44310cff44321dcf44311edf;
assign testcases[88] = 512'h10000fef10000fff963109df92100dff60100eff70100aef70421bbf70311bbf10100fff00000fff76541abf67431bcf56310aef664109ef57431cbf57411cbf;
assign testcases[89] = 512'h10010fef10000fffa73107dfa2100cff60100eff801109ef80421abf80421abf10110fff10000fff876429af78531abf66410aef775108ef69541baf68512bbf;
assign testcases[90] = 512'h00000fff10000fff41000fff50000fff20000fff30000fff30000fef30000fef00000fff00000fff21000fef21000fff21000fff21000fff21000fef21000fef;
assign testcases[91] = 512'h10000fef10000fff63100eff61000fff30000fff40000eff50210edf50100edf00000fff00000fff43211eef33210eef33200eff33200dff33210edf33201fdf;
assign testcases[92] = 512'h10000fef10000fff74200cef71000eff40100fff50100cff60210ddf60211ddf10000fff00000fff54321ddf44321ddf44210dff44310cff45321ddf45311edf;
assign testcases[93] = 512'h10000fef10000fff86210adf91100eff50100fff60100bff70311ccf70311ccf10000fff00000fff65431bcf56431ccf55310cff55410aef56431dcf56411dcf;
assign testcases[94] = 512'h10000fef10000fff973109df92100dff60100eff70100aef70421bbf70311bbf10000fff00000fff76541abf67431bbf66310bef664109ef68431cbf57412cbf;
assign testcases[95] = 512'h10010fef10000fffa83107cfa2100cff70100eff801109ef80421abf80421abf10110fff10000fff876429af78541abf67410aef775108ef69541bbf68512baf;
assign testcases[96] = 512'h00000fff10000fff52000fff50000fff20000fff30000fff30000fef40000fef00000fff00000fff21000fef21000fff21000fff21000fff22000fef22000fef;
assign testcases[97] = 512'h10000fef10000fff63100eff61000fff30000fff40100eff50210edf50100edf00000fff00000fff43211eef43210eef33200eff33200dff33210edf33200edf;
assign testcases[98] = 512'h10000fef10000fff74200cef71000eff40100fff50100cff60310dcf60211ddf10000fff00000fff54431cdf55321ddf44310dff44310cff45321dcf45311dcf;
assign testcases[99] = 512'h10000fef10000fff86210adf82100eff50100fff60100bff70311ccf70311ccf10000fff00000fff65431bcf56431ccf55310cff55410bef56431dcf56411dcf;
assign testcases[100] = 512'h10000fef10000fff973109dfa2100dff60100eff70100aff70421bbf80311bcf10110fff10000fff86542abf67431bcf66310bff664109ef68431cbf57412cbf;
assign testcases[101] = 512'h10010fef10100fffa83107cfa2100cff70110eff801109ef80421abf80421abf10110fff10000fff976428af79541abf67410aef775108ef69541bbf69512baf;
assign testcases[102] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff30000fef40000fef00000fff00000fff21000fef21000fff21000fff21000fff21000fef21000fef;
assign testcases[103] = 512'h10000fef10000fff63100eff61000fff30000fff40100eff50210edf50100edf00000fff00000fff42211edf43210eef32200eff33200dff33210edf33200edf;
assign testcases[104] = 512'h10000fef10000fff74200cef71000eff40100fff50100cff60310dcf60211dcf10000fff00000fff53431ccf54321ddf44310dff54310cff44321dcf44311dcf;
assign testcases[105] = 512'h10000fef10000fff95210adf91100eff50100fff60100bff70311ccf70311ccf10000fff00000fff64541bbf65431ccf55310bff65410aef56431ccf55411dcf;
assign testcases[106] = 512'h10000fef10000fffa73108dfa2100dff60100eff70100aef80421bbf80421bbf10100fff00000fff866429af77541abf66410aef665109ef67541bbf67512cbf;
assign testcases[107] = 512'h10010fef10100fffb83107cfb2100cff70100eff801109ef80421aaf80421abf10110fff10000fff976528af785419bf674109ef775108ef69541baf69512baf;
assign testcases[108] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff40000fef40000fef00000fff00000fff21000fef21000fef21000fff21000fff21000fef21000fef;
assign testcases[109] = 512'h10000fef10000fff63100eef61000fff30100fff40100eff50210edf50210edf00000fff00000fff43221edf43210eef33200eff33200dff33210edf33201edf;
assign testcases[110] = 512'h10000fef10000fff84200cef81100eff40100fff50100cff60311dcf60311dcf10000fff00000fff64431ccf55321ddf44310dff54310cff45321dcf45311dcf;
assign testcases[111] = 512'h10000fef10000fff96210adf92100eff50100fff60100bff70311ccf70311ccf10000fff00000fff75541bbf66431ccf55310bff65410aef56431ccf56411ccf;
assign testcases[112] = 512'h10000fef10000fffa83109dfa2100dff60100eff70100aff70411bbf70411bbf10100fff10000fff87642abf68531bcf66410bef665109ef6a531cbf59511cbf;
assign testcases[113] = 512'h10010fef10000fffb83107cfb2100cff70110eff801108ef80421aaf80421aaf10110fff10000fff9765289f78541abf664109ef775108ef69541baf69512baf;
assign testcases[114] = 512'h00000fff10000fff52000fff50000fff20000fff30000fff30000fef40000fef00000fff00000fff31000fef21000fef21000fff21000fff22000fef22000fef;
assign testcases[115] = 512'h10000fef10000fff63100eff61000fff30000fff40100eff50210edf50100edf00000fff00000fff43221edf43210eef33200eff33200dff34210edf33201edf;
assign testcases[116] = 512'h10000fef10000fff74200cef81100eff40100fff50100cff60310dcf60211dcf10000fff00000fff54431ccf55321ddf44310dff44310cff45321dcf45311dcf;
assign testcases[117] = 512'h10000fef10000fff96310adf92100eff50100fff60100bff70411ccf70311ccf10000fff00000fff75541bbf66431ccf55310cff55410aef57431ccf56411dcf;
assign testcases[118] = 512'h10000fef10000fffa73108dfa2100dff60100eff70100aef70421bbf70311bbf10110fff10000fff866429af67541bbf66410aef664109ef68531bbf58512cbf;
assign testcases[119] = 512'h10010fef10100fffb83107dfb2100cff60110eff801109ef80421abf80421abf10110fff10000fff976528af78541abf67410aef775108ef69541baf69512baf;
assign testcases[120] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff30000fef40000fef00000fff00000fff21000fef21000fff21000fff21000fff22000fef22000fef;
assign testcases[121] = 512'h10000fef10000fff63100eff61000fff30000fff40000eff50210edf50100edf00000fff00000fff42211eef43210eef33200eff33200eff33210fdf33200fdf;
assign testcases[122] = 512'h10000fef10000fff74200cef71100eff40100fff50100cff60310ddf60211ddf10000fff00000fff53431ccf54321ddf44310dff44310cff45321dcf44311edf;
assign testcases[123] = 512'h10000fef10000fff85210adf81100eff50100fff60100bff60311ccf60311ccf10000fff10000fff65541bbf55431ccf55310cff55410bef56431ccf56411dcf;
assign testcases[124] = 512'h10000fef10000fff963109df92100dff60100eff70100aef70421bbf70311bbf10110fff10000fff76542abf67441bcf56310bef66410aef58431cbf57411cbf;
assign testcases[125] = 512'h10010fef10100fffb73107cfa2100cff60100eff701009ef80421abf80421abf10110fff10000fff966528af78541abf66410aef775108ef69541baf68512bbf;
assign testcases[126] = 512'h10000fef10000fff52100eff61000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef22100fff32100eff23110fef23100fef;
assign testcases[127] = 512'h10000fef10000fff74100def71000fff40100fff50100dff50210edf50210edf10000fff00000fff54321ddf44220edf33200dff43300dff35210edf35201edf;
assign testcases[128] = 512'h10000fef10000fff85200bef81100eff50100fff60100cff60311dcf60311dcf10000fff00000fff65531ccf55431ccf44310cff54410bff46321dcf46311dcf;
assign testcases[129] = 512'h10000fef10000fff962109df92100dff50100fff60100bff70311ccf70311ccf10000fff10000fff76542abf67431bcf55310bff65410aef57431ccf57411ccf;
assign testcases[130] = 512'h10010fef10100fffa83108dfa2100dff60100eff70100aef80421bbf80311bbf10110fff10000fff876429af78541abf66310aef664109ef69531bbf68512bbf;
assign testcases[131] = 512'h10000fef10000fff52100eff61000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef22100fff32100eff23110fef23100fef;
assign testcases[132] = 512'h10000fef10000fff74100def71000fff40100fff40100dff50210edf50210edf00000fff00000fff53321ddf44220edf33200eff43310dff35220edf34201edf;
assign testcases[133] = 512'h10000fef10000fff85200bef81100eff50100fff50100cff60311dcf60311dcf10000fff00000fff65431ccf56331cdf45310cff55310bff46321dcf46311dcf;
assign testcases[134] = 512'h10000fef10000fff973109df92100dff50100fff60100bff70311bbf70311cbf10100fff00000fff76541abf67431bcf55310bef66410aef58431cbf57411cbf;
assign testcases[135] = 512'h10000fef10100fffa83108dfa2100dff60100eff70100aef80421bbf80411bbf10110fff10000fff876529af78541abf66410aef664109ef69541bbf68512bbf;
assign testcases[136] = 512'h10000fef10000fff63100eff61000fff30000fff30000eff40100fef40100fef00000fff00000fff32210fef33110fef22100fff32100eff33110fef33100fef;
assign testcases[137] = 512'h10000fef10000fff74200def71000fff40100fff50100dff50210edf50210edf10000fff00000fff53321ddf44321ddf33200dff43310dff44221edf44201edf;
assign testcases[138] = 512'h10000fef10000fff85200bef81100eff50100fff60100cff60311ccf60311ccf10000fff00000fff65531bcf55431ccf44310cff55410bff46431dcf46411dcf;
assign testcases[139] = 512'h10000fef10000fff963109df92100dff60100fff70100aff70421bbf70311bbf10100fff10000fff76642abf67431bcf55310bff66410aef58431cbf57411cbf;
assign testcases[140] = 512'h10000fef10100fffa73107dfa2100cff60100eff801109ef80421abf80421abf10110fff10000fff967528af77541abf66410aef765108ef68541bbf68512baf;
assign testcases[141] = 512'h10010fef10100fffb93106cfb2100cff70110eff901108ef904219af904219af10110fff10110fffa875279f895519af774109ef875107ef7b541aaf7a512aaf;
assign testcases[142] = 512'h10010fef10100fffb83106cfb2100cff70110eff801108ef905219af904219af10110fff10010fffa875279f895519af774109ef875207ef7a541aaf79512aaf;
assign testcases[143] = 512'h10010fef10100fffb93106cfb2100cff70110eff801108ef905219af904219af10110fff10000fffa875279f895519af774109ef775107ef7a541aaf69512aaf;
assign testcases[144] = 512'h10000fef10000fff52100eff61000fff30000fff30000eff40100fef40100fef00000fff00000fff32210fef32110fef22100fff32200eff22110fef22100fef;
assign testcases[145] = 512'h10000fef10000fff73100def71000fff40100fff50100dff50210edf50210edf10000fff00000fff53321ddf43221edf33200dff43310dff34220edf33201edf;
assign testcases[146] = 512'h10000fef10000fff84200bef81100eff50100fff60100cff60311ccf60311ccf10000fff00000fff64531bcf54431ccf44310cff54410bff45431dcf45411dcf;
assign testcases[147] = 512'h10000fef10000fff953109df91100dff50100fff60100bef70411bbf70311cbf10100fff10000fff75542abf66431bcf55310bef65410aef57431cbf56411cbf;
assign testcases[148] = 512'h10000fef10100fffa73108dfa2100dff60100eff701109ef80421abf80421abf10110fff10000fff866529af77541abf66410aef765109ef68541baf67512bbf;
assign testcases[149] = 512'h10010fef10100fffb83106cfb2100cff70110eff801108ef904219af804219af10110fff10010fff9775279f885419af774109ef875107ef79541aaf79512baf;
assign testcases[150] = 512'h10000fef10000fff62100eff61000fff30000fff30000eff40100fef40100fef00000fff00000fff32210eef32110fef22100fff32200eff22110fef32100fef;
assign testcases[151] = 512'h10000fef10000fff74200cef71000eff40100fff50100dff50210ddf50211ddf00000fff00000fff53431ddf44321ddf43210dff43310cff44321edf44311edf;
assign testcases[152] = 512'h10000fef10000fff85210aef91100eff50100fff60100bff60311ccf60311ccf10000fff00000fff74541bcf55431ccf54310cff55410bef56431dcf56411dcf;
assign testcases[153] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff40000fef40000fef00000fff00000fff31000fef21000fef21000fff21000fff22000fef21000fef;
assign testcases[154] = 512'h10000fef10000fff63100def71000fff30100fff40100eff50210edf50110edf00000fff00000fff43321edf43210eef33200eff33200dff33210edf33201edf;
assign testcases[155] = 512'h10000fef10000fff84200bef81100eff40100fff50100cff60311dcf60311dcf10000fff00000fff64431ccf55331ddf44310dff54310cff45321dcf45311dcf;
assign testcases[156] = 512'h10010fef10100fffc94105cfb2100cff70110eff901107ef905219af904219af10110fff10000fffa886278f8965189f774108ef875206ef7a651aaf79612aaf;
assign testcases[157] = 512'h10010fef10100fffc94105cfc2100cff70110eff901108ef905219af904219af10110fff10010fffa876279f896519af774109ef875207ef7a641aaf79612aaf;
assign testcases[158] = 512'h00000fff10000fff52100fff61000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef22100fff32100eff23100fef23100fef;
assign testcases[159] = 512'h10000fef10000fff63100eff61000fff30000fff40000eff50100edf50100edf00000fff00000fff42211eef43210eef32200eff32200dff33210fdf33200fdf;
assign testcases[160] = 512'h00000fff10000fff52100fff60000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef32110fef22100fff32100eff22100fef22100fef;
assign testcases[161] = 512'h10000fef10000fff63100eff61000fff30000fff40000eff50110edf50100edf00000fff00000fff42221eef43210eef32200eff32200eff33210fdf33201fdf;
assign testcases[162] = 512'h00000fff10000fff52100fff61000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef22100fff32100eff22100fef22100fef;
assign testcases[163] = 512'h10000fef10000fff63100eff61000fff30000fff40000eff50110edf50100edf00000fff00000fff42211eef43210eef32200eff32200eff33210fdf33200fdf;
assign testcases[164] = 512'h10000fef10000fff52100fff51000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef22100fff22100fff23110fef23100fef;
assign testcases[165] = 512'h10000fef10000fff63100eff61000fff30000fff40000eff50100edf50100edf00000fff00000fff42210eef43210eef32100eff33200eff33110fdf33100fdf;
assign testcases[166] = 512'h10000fef10000fff52100fff61000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef32110fef22100fff32100eff22100fef22100fef;
assign testcases[167] = 512'h10000fef10000fff62100eff61000fff30000fff40000eff50210edf50100edf00000fff00000fff42221eef33210eef32200eff32200eff33210fdf33200fdf;
assign testcases[168] = 512'h10000fef10000fff52000fff50000fff20000fff30000fff40100fef40100fef00000fff00000fff31110fef32110fef22100fff22100fff22100fef22100fef;
assign testcases[169] = 512'h10000fef10000fff63100eff61000fff30000fff40000eff50100edf50100edf00000fff00000fff42211eef33210eef32100eff33200eff33210fdf33200fdf;
assign testcases[170] = 512'h10000fef10000fff52000fff61000fff30000fff30000fff40100fef40000fef00000fff00000fff32100fef32100fef22100fff32100eff22100fef22100fef;
assign testcases[171] = 512'h10000fef10000fff63100eff61000fff30000fff40000eff50210edf50100edf00000fff00000fff42211eef43210eef32200eff33200dff33210fdf33200fdf;
assign testcases[172] = 512'h10000fff10000fff64000fff61000fff30000fff40000fff40000fef50000fef00000fff00000fff43000fff44000fef33000fff33000fff34000fef34000fef;
assign testcases[173] = 512'h10000fef10000fff61000fff70000fff40000fff50000eff40100fef50000fef00000fff00000fff41100fef42100fef43100eff43100eff31100fef31100fef;
assign testcases[174] = 512'h10000fef10000fff61100fff70000fff50000fff60000cff50100fef50100fef00000fff00000fff41211fef52210fef53200dff53200cff31110fef31100fef;
assign testcases[175] = 512'h10000fef10000fff61100fff70000fff60100fff70100bff50100fef50100fef10000fff00000fff51221fef52221eef64200cff64300bff31210fef31200fef;
assign testcases[176] = 512'h10000fef10000fff61100fff70000fff70100fff80100aff50100fef50100fef10000fff00000fff51321fef63310eef64300bff74300aff31210fef41200fef;
assign testcases[177] = 512'h10000fef10000fff61100eff70000fff70100eff901009ff50200fef50200fef10000fff00000fff51321eef63421eef75310aef744109ef31210fef41201fef;
assign testcases[178] = 512'h10000fef10000fff61100eff80100fff80100eff901009ff50210fef50210fef10000fff00000fff51421eef63421eef75410aef744109ef41210fef41301fef;
assign testcases[179] = 512'h10000fef10000fff71200eff81100fff80100effa01008ef50210fef50210fef10000fff10000fff52432eef63432edf754109ef855108ef42321fdf42301fdf;
assign testcases[180] = 512'h10000fef10000fff72200eff81100fff90100effb01007ef50210fef60210fdf10000fff10000fef62421eef74421ddf864108ef965107ef42320fdf42301fdf;
assign testcases[181] = 512'h10000fef10000fff72200eff81100fffa0100dffc02006ef50210fef60211edf10110fff10100fef62531edf73531ddf965107ef966106ef42321fdf42311fdf;
assign testcases[182] = 512'h10000fef10100fff72200eff81100fffb0200dffd02104ef50310edf60311edf10110fff10110fef62641edf73641ddfa76106efa77105ef42431edf42411edf;
assign testcases[183] = 512'h10000fef10100fff72310def91100fffc0210dffe02103ef60311edf60311edf10110fff10110fef62642ddf74751ddfb77105efb78204ef42431edf42412edf;
assign testcases[184] = 512'h10000fef10100fff85310def92100fffc1200dffe02003ef60311edf60311edf10110fff10110fef65642ddf79751ddfbc6105efbb7104df55431edf55411edf;
assign testcases[185] = 512'h10110fef10100fff82310def91100effc0210cffe02102df60311edf60311edf10111fef10111fef62752ddf74862ccfb98104dfb89203df52531edf52512edf;
assign testcases[186] = 512'h10110fef10110fff82310cef91100effc0310cfff03101df60411edf60411edf10111fef10111fef62762ddf84962ccfc99203dfc9a202df52541edf52512edf;
assign testcases[187] = 512'h00000fff10000fff51000fff60000fff30000fff30000fff40000fef40000fef00000fff00000fff31000fff31000fff21000fff31000fff21000fef21000fef;
assign testcases[188] = 512'h00000fff10000fff61000fff60000fff40000fff50000eff40100fef40100fef00000fff00000fff41110fef42100fef32100eff42100eff31100fef31100fef;
assign testcases[189] = 512'h00000fef10000fff61100fff70000fff50000fff60000dff40100fef50100fef00000fff00000fff41210fef52210fef43100dff53200dff31110fef31100fef;
assign testcases[190] = 512'h10000fef10000fff61100fff71000fff60100fff70100bff50100fef50100fef00000fff00000fff52311fef53310eef64200bff64310bff32211fef32201fef;
assign testcases[191] = 512'h10000fef10000fff61100fff71000fff60100fff80100aff50100fef50100fef00000fff00000fff42311fef53320eef65200bff65300aef32210fef32200fef;
assign testcases[192] = 512'h10000fef10000fff62100eff71000fff70100eff801009ef50200fef50200fef10000fff00000fef52321eef63321edf66310aef754109ef32210fef32201fef;
assign testcases[193] = 512'h10000fef10000fff62100eff71100fff70100eff901009ef50210fef50210fef10000fff00000fff52421eef63421eef76310aef754109ef32210fef42201fef;
assign testcases[194] = 512'h00000fef10000fff61100fff70000fff50000fff60100cff40100fef50100fef00000fff00000fff41210fef53210fef44200dff53200cff31110fef31100fef;
assign testcases[195] = 512'h10000fef10000fff72200eff81100fff80100effa01008ef50210fef50210fef10000fff10000fff52421eef64421edf874109ef864108ef42321fdf42301fdf;
assign testcases[196] = 512'h10000fef10000fff72200eff81100fff90100effb01007ef50210fef50211fdf10110fff10000fef52431eef64531ddf874108ef875107ef42321fdf42312fdf;
assign testcases[197] = 512'h10000fef10000fff72200eff81100fffa0200dffc02005ef50310edf60311edf10110fff10110fef62541edf74641ddf985107ef976106ef42321edf42411edf;
assign testcases[198] = 512'h10000fef10100fff72210def81100fffb0200dffd02104ef50311edf60311edf10110fff10110fef62642ddf74751ddfa86106efa87105ef42431edf42411edf;
assign testcases[199] = 512'h10000fef10100fff82310def91100fffb0210dffe02103ef60311edf60311edf10110fff10110fef62652ddf74751cdfb97105efb88204ef42431edf42411edf;
assign testcases[200] = 512'h10110fef10110fff82310def91100effc0210dffe02102df60311edf60311edf10111fef10111fef63764ddf75863ccfba8204dfb99203df42551edf53512edf;
assign testcases[201] = 512'h10110fef10110fff82310cef91100effc0210cfff03102df60421edf60411edf10111fef10111fef63762ddf85962ccfca9204dfc99202df53541edf53512edf;
assign testcases[202] = 512'h00000fff10000fff51000fff60000fff30000fff30000fff40000fef40000fef00000fff00000fff31000fef31000fef21000fff21000fff21000fef21000fef;
assign testcases[203] = 512'h00000fff10000fff61000fff60000fff40000fff40000eff40100fef40100fef00000fff00000fff41110fef42100fef32100eff32100eff31100fef31100fef;
assign testcases[204] = 512'h10000fef10000fff61100fff71000fff60100fff70100cff40100fef50100fef00000fff00000fff42210fef53210eef54200cff54200cff31110fef32100fef;
assign testcases[205] = 512'h10000fef10000fff61100fff71000fff60100fff80100bff50100fef50100fef00000fff00000fff52321fef63310eef64200bff64300bff31210fef32200fef;
assign testcases[206] = 512'h10000fef10000fff61100fff71000fff70100eff90100aff50200fef50200fef10000fff00000fff52321fef63321eef75310aff75410aef31210fef42201fef;
assign testcases[207] = 512'h10000fef10000fff72100eff81100fff80100eff901009ef50210fef50210fef10000fff00000fff52421eef63421eef75410aef754109ef42210fef42301fef;
assign testcases[208] = 512'h10000fef10000fff72200eff81100fff80100effa01008ef50210fef50211fef10011fff00001fff52432eef63432edf864109ef855108ef42321fdf42311fdf;
assign testcases[209] = 512'h10000fef10000fff72200eff81100fff90100effb01006ef50210fef50210fef10000fff10000fef52431edf64531ddf864108ef865107ef42321fdf42311fdf;
assign testcases[210] = 512'h10000fef10000fff72200eff81100fffa0100dffc02006ef50210fef60211edf10110fff10000fef62531eef74531ddf975107ef966107ef42321fdf42311fdf;
assign testcases[211] = 512'h10000fef10100fff72200def81100fffb0200dffd02104ef50310edf60311edf10110fff10110fef62641edf74641ddfa86106efa77105ef42431edf42411edf;
assign testcases[212] = 512'h10000fef10100fff82310def91100fffc0210dffe02103ef60311edf60311edf10110fff10110fef62642ddf74751ddfb87105efb78104ef42431edf42411edf;
assign testcases[213] = 512'h10110fef10100fff82310def91100effc0210cfff02102ef60311edf60311edf10110fff10111fef62752ddf74851cdfb98204efb89203df42431edf52512edf;
assign testcases[214] = 512'h10110fef10100fff82310def91100effc0210cfff02102df60311edf60311edf10110fef10111fef62642ddf75751ddfba7104dfb98103df42431edf42411edf;
assign testcases[215] = 512'h10110fef10100fff72310def81100effc0210cffe02101df50311edf60311edf10111fef10111fee62652ddf74751dcfb97104dfb88103ef42431edf42411edf;
assign testcases[216] = 512'h10000fef10000fff61100fff70000fff50000fff60000dff40100fef40100fef00000fff00000fff41110fef52110fef43100dff43100dff31100fef31101fef;
assign testcases[217] = 512'h00000fff10000fff51000fff60000fff30000fff30000fff40000fef40000fef00000fff00000fff31000fff31000fef21000fff31000fff21000fef21000fef;
assign testcases[218] = 512'h00000fff10000fff51000fff60000fff40000fff50000eff40000fef40000fef00000fff00000fff41100fef42100fef32100eff42100eff31100fef31100fef;
assign testcases[219] = 512'h10000fef10000fff61100fff70000fff50000fff60000dff40100fef40100fef00000fff00000fff41210fef52210fef43100dff43200dff31100fef31100fef;
assign testcases[220] = 512'h10000fef10000fff61100fff70000fff60100fff70100cff40100fef50100fef00000fff00000fff41210fef52210fef54200cff54200cff31110fef31100fef;
assign testcases[221] = 512'h10000fef10000fff61100fff70000fff60100fff70100bff40100fef50100fef00000fff00000fff41211fef53310eef64200cff64300bff31210fef31200fef;
assign testcases[222] = 512'h10000fef10000fff61100fff70000fff70100eff80100aff50100fef50100fef10000fff00000fff51321fef53321eef65300bff65310aff31210fef31201fef;
assign testcases[223] = 512'h10000fef10000fff61100eff71000fff80100eff901009ef50200fef50200fef10000fff00000fff52321fef63421eef75310aef75410aef31210fef32201fef;
assign testcases[224] = 512'h10000fef10000fff61100eff71100fff80100effa01008ef50210fef50210fef10000fff10000fff52421eef63421eef764109ef754109ef31220fef42301fef;
assign testcases[225] = 512'h10000fef10000fff72200eff81100fff90100effb01007ef50210fef50211fef10011fff10001fef52431eef63532edf864108ef865108ef42321fdf42311fdf;
assign testcases[226] = 512'h10000fef10000fff72200eff81100fff90100effb01007ef50210fef50210fdf10000fff10000fef52421eef64421edf873108ef874108ef42210fdf42201fdf;
assign testcases[227] = 512'h10000fef10100fff72200eff81100fffa0100dffc02005ef50210fdf50211edf10110fff10110fef52531eef64541ddf975107ef976106ef42321fdf42311fdf;
assign testcases[228] = 512'h10000fef10100fff72200eef81100fffb0200dffd02104ef50310edf60311edf10110fff10110fef52541edf74641ddfa86106efa77105ef42331edf42411edf;
assign testcases[229] = 512'h10110fef10100fff72310def81100fffc0210cffe02102ef50311edf60311edf10110fff10110fef62652edf74761ddfb97105efa87104ef42431edf42411edf;
assign testcases[230] = 512'h10110fef10100fff72310def91100fffc0210cfff02102df50311edf60311edf10110fef10111fef62652ddf74862ddfb97104dfb88203df42431edf42512edf;
assign testcases[231] = 512'h10110fef10110fff82310def91100effd0310cfff03101df60311edf60311edf10111fef10111fef62752ddf74862ccfc98204dfb99203df42541edf42512edf;
assign testcases[232] = 512'h00000fff10000fff51000fff60000fff30000fff40000fff40000fef40000fef00000fff00000fff31000fff31000fff32000fff32000fff21000fef21000fef;
assign testcases[233] = 512'h00000fff10000fff51000fff60000fff40000fff50000eff40000fef40000fef00000fff00000fff41100fef42100fef32100eff42100eff31100fef31100fef;
assign testcases[234] = 512'h10000fef10000fff61100fff60000fff50000fff60000dff40100fef40100fef00000fff00000fff41110fef52210fef43100dff53200dff31100fef31100fef;
assign testcases[235] = 512'h10000fef10000fff61100fff70000fff60100fff70100cff40100fef50100fef00000fff00000fff41210fef52210fef54200cff53200cff31110fef31100fef;
assign testcases[236] = 512'h10000fef10000fff61100fff70000fff70100fff80100bff40100fef50100fef00000fff00000fff41211fef52320eef64310bff64310bff31210fef31201fef;
assign testcases[237] = 512'h10000fef10000fff61100fff70000fff70100eff80100aff50100fef50100fef10000fff00000fff51321fef53321eef64310bff74410aff31210fef31201fef;
assign testcases[238] = 512'h10000fef10000fff61100fff70000fff80100eff901009ef50200fef50200fef10000fff00000fff51321fef63421edf75310aef754109ef31210fef31201fef;
assign testcases[239] = 512'h10000fef10000fff61100eff81100fff90100effa01007ef50210fef50211fef10010fff10001fef52422eef63431edf854109ef855108ef41220fef42311fef;
assign testcases[240] = 512'h10000fef10000fff71200eff81100fff90100effb01007ef50210fef50210fef10000fff10000fff52431eef63531eef864108ef865108ef42321fdf42311fdf;
assign testcases[241] = 512'h10000fef10000fff72200eff81100fffa0100dffc02006ef50210fef50210fef10110fff10000fef52431eef63531edf965107ef966107ef42321fdf42311fdf;
assign testcases[242] = 512'h10000fef10100fff72200eff81100fffb0200dffd02004ef50210fdf50211edf10110fff10110fef52541edf73641ddfa76106efa66106ef42321fdf42411fdf;
assign testcases[243] = 512'h10000fef10100fff72210def81100fffc0210cffe02102ef50311edf60311edf10110fff10110fef62642edf74751ddfb87105efa77104ef42431edf42411edf;
assign testcases[244] = 512'h10110fef10100fff72310def91100fffd0210cfff02101df50311edf60311edf10110fff10110fef62652ddf74751ddfb87104dfb78204ef42431edf42411edf;
assign testcases[245] = 512'h10110fef10100fff82310def91100effd0210cfff03100df60311edf60311edf10111fef10111fef62752ddf74862cdfc98203dfc89202df42441edf42512edf;
assign testcases[246] = 512'h10110fef10110fff82310def91100effe0310cfff03100df60311edf60411edf10111fef10111fef62762ddf84972ccfc99203dfc8a202df42541edf52512edf;
assign testcases[247] = 512'h00000fef10000fff40000def40000eff20000cff200000df30000edf30000edf00000fef00000fef20000ddf20000cdf101003df201002df10000edf10000edf;
assign testcases[248] = 512'h30220edf30310def62100eff61000fff50100fff60100bff50210edf50211edf31331def31332ddf42321eef43321eef65510bff65510bff32321edf32311edf;
assign testcases[249] = 512'h40441ccf50420cef74200cef71000eff80110eff901108ef60311ccf60311ccf42442cdf52553bce53331ddf54321ddf875208ef876207ef44331dcf44311dcf;
assign testcases[250] = 512'h20220eef20210eff52100fff51000fff40100fff50100dff40110fef40100fef21221eef21221eef32210fef32110fef44310dff43310cff32110fef32201fef;
assign testcases[251] = 512'h50562fee50641fff84210cef91100fffa0210effb0210bff80423dcf80424dcf52664fef62776fee74554ddf75553ddfa9831befa8941aef65552dcf65622dcf;
assign testcases[252] = 512'h50561bbe50641bde95210ade91100effa0210dffb02106ef80521bad80421bbe52663ace627749bd74542bbe75541bbfa98317efa89316ef75642bae75612bae;
assign testcases[253] = 512'h00000fef10000fff51100eff60000fff30100fff40100dff40210edf40211edf00000fff00000fff31321eef31221eef32210eff32310dff31221edf31211edf;
assign testcases[254] = 512'h10000fef10100fffb65107dfb2110cff80210eff902109ef90732abf90632abf10110fff10000fff869839bf968729bf776209ef868208ef76772bbf75823bbf;
assign testcases[255] = 512'h10000fef10100fffa64109dfa2110dff70210eff80210aff80632bcf80632bcf10100fff10000fff85873abf76762abf77620aef76620aef66772ccf65723ccf;
assign testcases[256] = 512'h10000fef10100fffa64109dfa2110dff70210eff802109ef80631bbf80632bbf10100fff10000fff85873abf77762abf76620aef76720aef66772cbf66723cbf;
assign testcases[257] = 512'h10000fef10000fff62100eff61000fff40100fff40100eff50210edf50210edf00000fff00000fff42321eef42220eef33210eff43210dff32220edf32201edf;
assign testcases[258] = 512'h10000fef10100fffa64108dfa2110dff70210eff802109ef80631bbf80532abf10100fff10000fff85873abf86762abf76620aef766209ef66772bbf65723bbf;
assign testcases[259] = 512'h10000fef10000fff63100eff61000fff40100fff40100dff50210edf50210edf00000fff00000fff42321eef43220eef33210eff43210dff32210edf32201edf;
assign testcases[260] = 512'h10000fef10100fffa64108cfa2100dff70210eff802109ef80631aad80532aae10000fff10000fff858739ad867629ae776209ef766208ef65762baf65723bae;
assign testcases[261] = 512'h10221fef10220fff833109df91100dff70210eff802108ef80621aaf70522aaf10231fff10221fff62762aaf63651abf758218ef758207ef63762baf63723baf;
assign testcases[262] = 512'h10000fef10100fff944108dfa1100dff70210eff802108ef80631abf80532abf10000fff00000fff73773abf74762abf766209ef766208ef64662bbf64623bbf;
assign testcases[263] = 512'h10000fef10000fffa44108dfa1100dff70210eff802108ef80631abf80532abf10000fff00000fff74873abf75762abf776209ef766208ef64662bbf64723bbf;
assign testcases[264] = 512'h10672fef10861eef72510def81210effa0310dffc03105ef50731edf60722dcf10794eef10785eef51a73ddf62b72ddfa7b206efa7c205ef31862ecf41823ecf;
assign testcases[265] = 512'h10110fef20210eff72310def81100effc0310cffd03102df50421edf60421edf10221eef10221eef51642ddf62751ddfb99204dfb8a203df31431ecf41411edf;
assign testcases[266] = 512'h10110fef10110fef72310def81100effc0210cffe03101df50421edf60421edf10221eef10221eee51642ddf62751dcfb99203dfb89202df31431edf41411edf;
assign testcases[267] = 512'h10110fef20110eff72310def91100effc0310cffe03102df60311edf60311ddf10111eef11111eef52542ddf63751ddfc98203dfc89203df42431ecf42411edf;
assign testcases[268] = 512'h10110fef10110fff72310def81100effc0210cffe03102df50311edf60411edf10111fef10211fef52542ddf63751ddfc98204dfb89203df42431edf42411edf;
assign testcases[269] = 512'h10111fef20111eef72310cef91110effc0311cffe03111df60423edf60424ddf11223eef11223eef52666ddf63786ccfc9a203dfc8b212df41431edf42412edf;
assign testcases[270] = 512'h10110fef10110fff72310def91100effc0310cffe03102df60312edf60421edf10121eef10112eef52543ddf63752ddfc99203dfc89203df42441edf42411edf;
assign testcases[271] = 512'h20110fef20110eff41000fff50000fff20000fff30000fff30000fef30000fef21110eef21111fef21000fff21000fff22100fff22100fff21000fef21000fef;
assign testcases[272] = 512'h30210ede30210def51000fff50000fff30000fff30000fff40100fef40000fef31221def31221ddf21100fef21100fef22100fff32100eff21100fef21100fef;
assign testcases[273] = 512'h30221ddf40320def52000fff50000fff30000fff40000eff40100fef40100fef41331ddf31332dde31110fef32110fef33200eff32200eff22110fef22100fef;
assign testcases[274] = 512'h40331dcf40420cef52000fff50000fff30000fff40000eff40100fef40100fef41442cdf41442cce31110fef32110fef33200eff33200eff22110fef22100fef;
assign testcases[275] = 512'h40441ccf50430bdf52100fff51000fff40100fff40100eff40100fef40100fef51442bdf41442bce32110fef32110fef33210eff43310dff22110fef32100fef;
assign testcases[276] = 512'h50551bbe60631adf52100eff61000fff40100fff50100dff50100edf50100edf51663acf52663abe32210fef33110fef44310dff44310cff33110fdf33201fdf;
assign testcases[277] = 512'h60661abe706419cf63100eff61000fff50100fff50100cff50210edf50100edf627739cf627749ae43211eef43210eef44310dff54310cff33210edf33201edf;
assign testcases[278] = 512'h60772aae707518ce63100def61000fff50100fff60100cff50210edf50210edf728838be728849ae43221edf44210edf55310cff55410bff34210edf44201edf;
assign testcases[279] = 512'h707729ae808518ce64100def71000fff50100fff60100bff60210ddf60210ddf828848be8288589e43221ddf44210edf55410cff65410bef44220edf44201ecf;
assign testcases[280] = 512'h707829ae808617ce74100def71000fff60100fff70100bff60210dcf60210dcf828947ae8289579e54221ddf44220ddf66310bef66410aef45220dcf45201dcf;
assign testcases[281] = 512'h8088289e909617be74100cef71000eff60100eff70110aef60210ccf60211dcf929a47ae8299579d54321ddf54320ddf66410aef66410aef45321dcf45311dcf;
assign testcases[282] = 512'h8099289d90a616be75200cef71000eff70100eff801109ef60310ccf60211ccf92aa46ae92aa578d54321ccf55320ccf67410aef765109ef55321ccf55311dcf;
assign testcases[283] = 512'h909a279da0a716be75200bef81000eff70100eff801109ef70310cbf70211ccf92ab56ae92aa668d54321ccf55321ccf774109ef775108ef56321cbf55311cbf;
assign testcases[284] = 512'h909b378da0a716ad85200bef81000eff70110eff801108ef70310bbf70211bbfa2ac669da2ac767c65321bcf56321bcf774109ef774108ef56321cbf56311cbf;
assign testcases[285] = 512'h90ab378da0b816be86200adf81000eff80110eff901107ef80310abf70311bbfa2bc559ea2ac768d65421bbf66321bbf884108ef875107ef66421baf66411baf;
assign testcases[286] = 512'h90ab37ffa0b816ff86200aff81000eff80110eff901107ff80310aff80311bffa2bc65ffa2bc76ff65321bff66321bff874108ff875107ff66321bff66411bff;
assign testcases[287] = 512'h909a279da0a716bd85200adf81000eff80110eff901108ef70310baf70311bafa2ab569da2aa668c65421bbf66321bbf774108ef875107ef66421baf56411baf;
assign testcases[288] = 512'h9099289d90a716be85200bef81000eff70100eff801108ef70310bbf70311bbf92ab56ae92aa678d64321ccf55321ccf774109ef775108ef56321cbf55411cbf;
assign testcases[289] = 512'h20110fef20110eff41000fff50000fff20000fff30000fff30000fef30000fef20110eef20111eef21000fff21000fff21100fff21100fff21000fef21000fef;
assign testcases[290] = 512'h20220ede30210def51000fff50000fff30000fff30000fff40000fef40000fef31221def31221dde21100fef21100fef32100fff32100eff21000fef21100fef;
assign testcases[291] = 512'h30221dde40320def52000fff50000fff30000fff40000eff40100fef40100fef41331dde31332dde31110fef31100fef32200eff32200eff22100fef22100fef;
assign testcases[292] = 512'h40331dce40420cde52000fff51000fff30100fff40100eff40100fef40100fef41442cdf41442cce32110fef32110fef33200eff43200dff22110fef22100fef;
assign testcases[293] = 512'h40441cce50430bdf52100fff51000fff40100fff40100dff40100fef40100fef51442bdf41442cce32110fef32110fef43210eff43310dff32110fef32100fef;
assign testcases[294] = 512'h50551bbe60631acf63100eff61000fff40100fff50100dff50100edf50100edf51663abf51563aad32210eef33210eef44310dff44310cff33210fdf33200edf;
assign testcases[295] = 512'h60561abe707419ce63100eff61000fff50100fff60100cff50210edf50200edf617739ce62674abe43211eef43210eef54310cff54410cff33210edf33201edf;
assign testcases[296] = 512'h60662aae707419ce63100def61000fff50100fff60100bff50210ddf50210edf727738be7277499d43211edf44210edf55310cff55410bff44210edf44201edf;
assign testcases[297] = 512'h7077299d808518be74100def71000fff60100fff70100bff60210dcf60210dcf828848ad7288589d53321ddf44210ddf65410bff65410aef44320dcf44301dcf;
assign testcases[298] = 512'h708829ae809518ce74100cef71000eff60100eff70100aef60310ccf60210dcf829947be8299589e54321ddf54320ddf66410aef65510aef45321dcf44311dcf;
assign testcases[299] = 512'h8088289d909616be74200cef71000eff60100eff80100aef60310ccf60210ccf9299469d8299577c54321ccf55320ddf66410aef765109ef55321dcf55311dcf;
assign testcases[300] = 512'h8098288d90a616bd75200bef81000eff70110eff801109ef70310cbf70311ccf92a9469d92a9577c54321ccf55320ccf76410aef765109ef55321cbf55311cbf;
assign testcases[301] = 512'h30110fef30100eef41000fff50000fff20000fff30000fff30000fef30000fef30110eef30111eef21000fff21000fff21000fff21000fff21000fef21000fef;
assign testcases[302] = 512'h40110dde50210cef51000fff50000fff30000fff30000fff40000fef40000fef50212cdf51212dde21000fef31000fff32000fff32100fff21000fef21000fef;
assign testcases[303] = 512'h50221cce60310bdf51000fff50000fff30000fff40000eff40000fef40000fef61321bcf61322bce31000fef31000fef32100eff32100eff21000fef21000fef;
assign testcases[304] = 512'h70331bbe80420ade52000fff50000fff40000fff40000eff40100fef40000fef71432ace71432abe31100fef32100fef43100eff43100eff32100fef32100fef;
assign testcases[305] = 512'h80543aae905309ce52000eff61000fff40000fff50000dff50100fef50100fef815529be815579ae32111fef32100fef43100eff43200dff32100fdf32100fdf;
assign testcases[306] = 512'h806519ae906318ce62000eff61000fff40000fff50000dff50100edf50100edf916537be9165389d42110eef42110eef44200dff43200dff32100edf32100edf;
assign testcases[307] = 512'h9065189ca06317be62100eef61000fff50000fff60000dff50100edf50100edfa16637ad9166378c42110edf42110edf54200dff53200cff42110edf42100edf;
assign testcases[308] = 512'h9076288da07417be63100eff61000fff50100fff60100cff50100edf50100edfa176379ea177478d42110eef43110eef54200dff54200cff42110edf42100edf;
assign testcases[309] = 512'ha087278db09516be73100def71000fff60100fff60100cff60200ddf60100ddfb19845aeb198568d53210ddf53210ddf54300cff64300bff43210ddf43200dcf;
assign testcases[310] = 512'hb099257cc0a514ad84100cef81000eff60100fff70100bff70210ccf70200ccfc1a9448dc1a9547d63211cdf54210cdf65310bff65310aff54210ccf53201ccf;
assign testcases[311] = 512'hc0ba355cd0b6139d84100bef81000eff70100eff80100aff70310bcf70210ccfd1bb537cd1bb645b63321ccf64310ccf75310aef75410aef54310ccf64301cbf;
assign testcases[312] = 512'he0cb334be0c7129d95200adf91000eff80100eff901009ef80310aaf80310abfe1cc627ce2cc725a74421bbf75321bbf864109ef864108ef75421baf75401baf;
assign testcases[313] = 512'hf0ee424af0e8119d952009df91100dff80100eff901008ef904109af90311abff1ee717cf2ee814a75421abf76421abf874108ef865108ef76521aaf75511aaf;
assign testcases[314] = 512'hf0ff4139f0f9208ca62008dfa2100dff80100effa01007efa04119af904119aff1ff705bf2ff9029855319bf865219bf985108ef975107ef865319af8651199f;
assign testcases[315] = 512'h30000fef30000eff41000fff50000fff20000fff30000fff30000fef30000fef30000eef31000fef21000fff21000fff21000fff21000fff21000fef21000fef;
assign testcases[316] = 512'h40110dde50210cef51000fff50000fff30000fff40000fff40000fef40000fef51211cdf51111dde31000fef31000fef32000fff32100fff21000fef21000fef;
assign testcases[317] = 512'h50221cce60310bdf51000fff50000fff30000fff40000eff40000fef40000fef61321bde61321bce31000fef31000fef32100eff32100eff21000fef31000fef;
assign testcases[318] = 512'h70331bbe80420ade52000fff60000fff40000fff50000eff50100fef50000fef71432ace71432abe31100fef32100fef43100eff43100eff32100fef32100fef;
assign testcases[319] = 512'h80441aae905219ce62000eff61000fff40000fff50000dff50100edf50100edf815438be815439ae42100eef42100eef43100dff43200dff32100fdf32100edf;
assign testcases[320] = 512'h905519ada06317ce62100eff61000fff50000fff60000dff50100edf50100edf916527be9165389d42110edf42110eef53200dff53200cff42110edf42100edf;
assign testcases[321] = 512'h9066289da07417be63100def71000fff50100fff60100cff60100ddf60100edfa17637aea176478d42110edf43110edf54200cff53200cff42110edf42100edf;
assign testcases[322] = 512'ha077278db08416be73100def71000fff50100fff60100cff60100ddf60100ddfb18736ada187468d52210ddf53210ddf54200cff64300bff43210ddf43200dcf;
assign testcases[323] = 512'hb098267cc0a515ad73100cef71000fff60100fff70100bff70200ccf60200dcfb1a9459db199557c53210dcf53210ddf64310bff64310bff53210dcf53200dcf;
assign testcases[324] = 512'hb0a9367dc0b615ae73100cef71000eff60100fff70100bff70210ccf70210ccfc1ba549dc1aa657d53311cdf53210ddf65310bff64410bff53310dcf53301dcf;
assign testcases[325] = 512'hd0bb346cd0c613ad84200bef81000eff70100eff80100aff80310bbf80210bcfd1cb538dd1cb736b63321bcf64320bcf75410aef754109ef64321bbf64301bbf;
assign testcases[326] = 512'he0cc324bf0d7129c952009df91000dff80100eff901008ef90310aaf80310aaff1dc627cf2cc725a74421abf75320abf864109ef864108ef75421aaf75411aaf;
assign testcases[327] = 512'hf0ff414bf0f8219ca52008dfa1100dff80100effa01008ef904119af904119aff1fe717cf1ff9149845319af855219af875108ef865107ef855319af855119af;
assign testcases[328] = 512'hf0ff400af0f9206ca63007cea1100cff90100dffa01006efa051189fa041189ff1ff704cf1ffa0098563189f8653189e975107ef975106ef8663199f8561199f;
assign testcases[329] = 512'h30110fef30100eff41000fff50000fff20000fff30000fff30000fef30000fef30110eef30111eee21000fff21000fff21000fff21000fff21000fef21000fef;
assign testcases[330] = 512'h40220dde50211cef51000fff50000fff30000fff40000fff40000fef40000fef50222cdf51223cde31000fef31000fef32100fff32100fff21000fef21000fef;
assign testcases[331] = 512'h50321cbe60310bde51000fff50000fff40000fff40000eff40000fef40000fef61321bce61322bbd31100fef31100fef32100eff42100eff31100fef31100fef;
assign testcases[332] = 512'h70431bbe804209ce62000eff60000fff40000fff50000eff50100eef50100fef714429ce71442abe31100fef32100fef43100eff42100dff32100fdf31100fdf;
assign testcases[333] = 512'h70541aae805308ce62100eff61000fff50000fff50000dff50100edf50100edf815428be815439ad42110eef42110eef53200dff53200dff42100edf42100edf;
assign testcases[334] = 512'h806519ad906318ce62100def71000fff50100fff60100cff60100ddf60100edf916537be9165389d42210edf42110edf53200cff53200cff42110edf42200edf;
assign testcases[335] = 512'h9076289da07417be72100def71000fff50100fff60100cff60200ddf60100ddfa17637aea176479d52210ddf52210ddf54200cff53300cff42210ddf42200ddf;
assign testcases[336] = 512'ha076278db07416be73100def71000fff60100fff70100cff60100ddf60100ddfb17636aea176468d52210ddf53210ddf64200cff64300bff53210dcf53200dcf;
assign testcases[337] = 512'hb098267cc09515ad83100cef81000eff60100fff70100bff70210ccf70200ccfc198459db198557c63311cdf63210cdf64310bff64410aff53310ccf53301ccf;
assign testcases[338] = 512'hc0aa346cd0b6139d93200aef81000eff70100eff801009ef80310bbf80310bbfd1ba538dd1ba646b63321bcf64321bcf75410aef744109ef64321bbf63301bbf;
assign testcases[339] = 512'hc0cb345cd0c7139d93200adf91100eff70100eff801009ef80410bbf80311bbfd1cc638dd1cc736c73421bcf64421bcf75410aef755109ef64421bbf63411bbf;
assign testcases[340] = 512'he0dc325af0d7129da42009dfa1100dff80100effa01008ef904109af90311aafe1dd627ce1dc724b84421abf85421abf864109ef855108ef85421aaf74411aaf;
assign testcases[341] = 512'hf0ee4139f0f8218cb53008dfa1100dff90100effa01007efa051189fa04119aff1fe717cf1ee914a946319af855319af975108ef966107ef8563199f8561199f;
assign testcases[342] = 512'hf0ff403af0f9208bb63106cfb1100cff90200dffb02006efb062179db051189ef1ff706bf1ffa039956318ae966318afa75107efa76106ef9673188d9571188d;
assign testcases[343] = 512'hf0ff4139f0f9208cb63106cfb1100cff90100dffb02006efb062179fb051179ff1ff706bf1ff9039956318af966317afa75107efa76106ef9673189f9571188f;
assign testcases[344] = 512'hf0ef614af0f8218cb53007dfa1100dff90100effa01007efa051189fa04118aff1efa16bf1ef913a956329af955318af975108ef975107ef9663199f8561299f;
assign testcases[345] = 512'hf0a9225bf0a6129da62009dfa2000dff80100effa01008efa03109af902109aff2a9427cf2a9625b85321abf873209bf973108ef874108ef87310aaf86301aaf;
assign testcases[346] = 512'he076235bf073139d971009df92000dff80100eff901009ef90210abf90200abff376328ce376336b76311abf77210abf872009ef873008ef78310abe77301aae;
assign testcases[347] = 512'hc0aa346cd0b614ad94200adf91000eff70100eff801009ef80310abf80310bbfd1ba538dd1aa646b73321bbf74320bbf75410aef754109ef74321bbf64301bbf;
assign testcases[348] = 512'hb098267dc09515ae83100bef81000eff70100fff80100aff70210ccf70210ccfc199448db199557c63311ccf63310ccf74310bff74410aff63310ccf63301ccf;
assign testcases[349] = 512'ha077279db08416be73100cef71000eff60100fff70100bff70200ccf70200dcfa18736ada187468d52210ddf53210ddf64300cff64300bff53210dcf53200dcf;
assign testcases[350] = 512'h9066189da07417be72100def71000fff60100fff70100cff60200ddf60100ddf917637ad9176478d52210ddf52210ddf64200cff63300bff52210ddf52200dcf;
assign testcases[351] = 512'h805519ae906318ce72100def71000fff50100fff60100cff60100ddf60100ddf916538be9165389d52210edf52110edf53200cff53200cff42210edf42200edf;
assign testcases[352] = 512'h70541aae805209ce62100eff61000fff50000fff60000dff60100edf60100edf815428be815439ae42110eef42110eef53200dff53200cff42110edf42100edf;
assign testcases[353] = 512'h60431bbe70420ade62000eff60000fff40000fff50000dff50100edf50100edf71432ace71432abe41110eef42100eef43100dff42200dff32100fdf31100edf;
assign testcases[354] = 512'h50321cce60310bde61000fff60000fff40000fff50000eff50100fdf50100fef61321bce61322bce31100fef31100fef42100eff42100eff31100fdf31100fdf;
assign testcases[355] = 512'h40210dce50210cde51000fff50000fff30000fff40000fff40000fef40000fef50221cdf40221dce31000fef31000fef32100fff32100eff21000fef31000fef;
assign testcases[356] = 512'h30110fef30100eff41000fff50000fff30000fff30000fff40000fef40000fef30110eef30111eef21000fff21000fff21000fff21000fff21000fef21000fef;
assign testcases[357] = 512'h30110fef30100eef51000fff50000fff30000fff30000fff40000fef40000fef30110eef30111eef21000fff21000fff21000fff21000fff21000fef21000fef;
assign testcases[358] = 512'h40110dde50210cef51000fff50000fff30000fff40000fff40000fef40000fef51211cdf51211dde31000fef31000fef32100fff32100eff21000fef31000fef;
assign testcases[359] = 512'h60221cce60310bde51000fff60000fff40000fff50000eff50000fef50000fef61321bce61321bce31100fef31100fef42100eff42100eff31100fef31100fef;
assign testcases[360] = 512'h70431bbe804209ce62000eff60000fff40000fff50000dff50100edf50100edf714329be71432aad41100eef42100eef43100dff42200dff32100fdf32100edf;
assign testcases[361] = 512'h805419ae905308ce62100eff71000fff50000fff60100dff60100edf60100edf815428be815439ad42110eef42110eef53200dff53200cff42110edf42100edf;
assign testcases[362] = 512'h8065189d906317be72100def71000fff50100fff60100cff60100ddf60100ddf916537ad9165388c52210ddf52210ddf53200cff53300cff42210edf42200edf;
assign testcases[363] = 512'h9076289da07417be73100def71000fff60100fff70100cff70200ddf60200ddfa17636aea176478d52210ddf53210ddf63300cff63300bff52210dcf52200dcf;
assign testcases[364] = 512'ha087278db08416be83100cef81000eff60100fff70100bff70210ccf70200ccfb18736ada187468d52211ddf53210ddf64310bff64310bff53210dcf53201dcf;
assign testcases[365] = 512'hb099267cc0a515ae83200bef81000eff70100eff80100aff80310bcf70210ccfc1a9459db1a9557c63321ccf63320ccf74410bff74410aff63320ccf63301cbf;
assign testcases[366] = 512'hc0ba356cc0b6149d94200aef91000eff70100eff80100aef80310bbf80310bbfc1ba547dc1ba645c73421bcf74321bcf75410aef745109ef64421bbf63411bbf;
assign testcases[367] = 512'hd0cc636be0c7339da42009dfa1100dff80100eff901009ef904119af90311abfe1ccc38cd1ccd36b83422abf74421abf855109ef855118ef74422aaf74513aaf;
assign testcases[368] = 512'he0dd325af0d8129da53008dfa1100dff90100effa01008efa05118afa04119afe1dd627ce1dd824b845319af855319bf965108ef966107ef855319af8451199f;
assign testcases[369] = 512'hf0ee4129f0f8217bb53106beb1100cff90100dffb02006efb051178db051178ef1fe715bf1ee812a9463188d9563188e975107ef966106ef9563188d9561188d;
assign testcases[370] = 512'hf0ff4138f0f9208cc63106cfc1100cffa0200dffb02006efc062168eb051179ff1ff706cf1ff904aa574179fa674179fa76106efa76106efa674178ea571278f;
assign testcases[371] = 512'h30331edf40320def52000fff51000fff40100fff40100dff40100fef40100fef41442def41332ddf32110fef33110fef44200dff44200dff33110fef33100fdf;
assign testcases[372] = 512'h40331dde50420cef51000fff50000fff30000fff40100eff40100fef40100fef51442cdf41442dce21110fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[373] = 512'h40341ddf50430cef52000fff50000fff30000fff40000eff40100fef40100fef51552cdf41442dde21100fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[374] = 512'h40441dde50530cde52000fff50000fff30000fff40000eff40100fef40100fef51552cde52542cce31100fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[375] = 512'h40441dde50530cef52000fff50000fff30000fff40100eff40100fef40100fef51552bdf52553cde31110fef32110fef33200eff43200dff22100fef22100fef;
assign testcases[376] = 512'h40441dde50531cde52000fff50000fff30100fff40100eff40100fef40100fef62552bde52553cde31110fef32110fef33210eff43200dff22100fef32100fef;
assign testcases[377] = 512'h40441dde50531cde52000fff50000fff40000fff40100eff40100fef40100fef62552bde52553cde31110fef32110fef44210dff43200dff22100fef32100fdf;
assign testcases[378] = 512'h40441ddf60531cef52000fff51000fff40100fff40100eff40100fef40100fef62552bdf52553cde32110fef32110fef44210dff43200dff22110fef32100fef;
assign testcases[379] = 512'h40451dce60631cde52000fff51000fff40100fff40100dff40100fdf40100fdf62663bce52563cce32110fef32110eef44210dff44310dff22110fdf32100fdf;
assign testcases[380] = 512'h20110fef30210eef41000fff40000fff20000fff30000fff30000fef30000fef31221eef21221eee21000fff21000fff22100fff22100fff21000fef21000fef;
assign testcases[381] = 512'h30331ede40320def41000fff50000fff30000fff30000fff40000fef40000fef41332ddf41332dde21100fff21100fff33200fff32200eff21000fef21100fef;
assign testcases[382] = 512'h30331edf40420def41000fff50000fff30000fff40000eff40100fef40000fef41442cdf41442dde21100fff32100fef33200eff33200eff21100fef22100fef;
assign testcases[383] = 512'h40331dde50420cef51000fff50000fff30000fff40000eff40100fef40100fef51442cde41442dde21100fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[384] = 512'h40341dde50430cef52000fff50000fff30000fff40000eff40100fef40100fef51552cdf41442dde31100fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[385] = 512'h40441dde50530cef52000fff50000fff30000fff40100eff40100fef40100fef52552cdf42553cde31110fef32110fef33210eff33200eff22110fef22100fef;
assign testcases[386] = 512'h40441ddf50531cef52000fff50000fff30100fff40100eff40100fef40100fef52552bdf52553cde31110fef32110fef33210eff43210eff22110fef32100fef;
assign testcases[387] = 512'h40441dde50531cde52000fff50000fff30100fff40100dff40100fdf40100fdf62562bde52553cce31110fef32110fef43210dff43310dff22110fdf32100fdf;
assign testcases[388] = 512'h40441dde50531cde52000fff51000fff40100fff40100eff40100fef40100fef62663bdf52553cde31110fef32110fef43210dff43310dff22110fef32100fdf;
assign testcases[389] = 512'h40451dde60531cee52100fff51000fff40100fff40100eff40100fef40100fef62663bde52553cde32110fef32110fef43210dff43310dff22110fef32100fdf;
assign testcases[390] = 512'h40564dde60641cee52100fff51000fff40100fff40100eff40101fef40100fef62673bde5267acde32111fef32111fef44210dff43310dff22110fdf32101fdf;
assign testcases[391] = 512'h50551ddf60641cef52100fff51000fff40100fff40100dff40100fef40100fef62663bdf52663cce32110fef32110fef44210dff43310dff22110fef32100fef;
assign testcases[392] = 512'h10110fef20100fff41000fff40000fff20000fff20000fff30000fef30000fef20110fff10110fef20000fff20000fff21000fff21100fff10000fef10000fef;
assign testcases[393] = 512'h20110fef30210eff41000fff40000fff20000fff30000fff30000fef30000fef31221eef21221eef21000fff21000fff22100fff22100fff21000fef21000fef;
assign testcases[394] = 512'h20220ede30210eef41000fff50000fff20000fff30000fff30000fef30000fef31321def31221ede21000fff21000fff22100fff22100fff21000fef21000fef;
assign testcases[395] = 512'h30221edf40320def41000fff50000fff30000fff30000fff30000fef30000fef41331ddf31332dde21000fff21000fff22100fff32100fff21000fef21000fef;
assign testcases[396] = 512'h30331ede40320def41000fff50000fff30000fff30000fff30000fef30000fef41442cdf41332dde21000fff21100fff32100fff32200fff21000fef21100fef;
assign testcases[397] = 512'h30331ede40420dee41000fff50000fff30000fff30000fff40100fef40000fef41442cdf41442dde21100fef22100fef33200eff32200eff21100fef22100fef;
assign testcases[398] = 512'h40331dde50430cef51000fff50000fff30000fff40000eff40100fef40100fef51442cde41442dde21100fef32100fef33200eff33200eff22100fef22100fef;
assign testcases[399] = 512'h40441dde50430cef52000fff50000fff30000fff40000eff40100fef40100fef51552cdf41442dde31110fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[400] = 512'h40441dce50530cde52000fff50000fff30000fff40100eff40100fef40100fef51552cde51553cce31110fef32110fef33200eff33200eff22110fef22100fef;
assign testcases[401] = 512'h40441dce50531cde52000fff50000fff30100fff40100eff40100fef40100fef51552bce52553cce31110fef32110fef33210eff43210eff22110fef32100fef;
assign testcases[402] = 512'h40441dce50531cde52000fff50000fff30100fff40100eff40100fef40100fef62552bde52553cce31110fef32110fef43210eff43200dff22110fef32100fef;
assign testcases[403] = 512'h40441dde60531cee52000fff51000fff40100fff40100eff40100fef40100fef63552bde53553cce32110fef33110fef44210eff43310dff23110fef33100fef;
assign testcases[404] = 512'h40441dce60531cde52100fff51000fff40100fff40100eff40100fef40100fef62652bde52553cce32110fef32110fef43210dff43310dff22110fef32100fdf;
assign testcases[405] = 512'h50451dde60531cee52000fff51000fff40100fff40100dff40100fdf40100fdf62652bde52553cde32110fef32110fef44210dff43210dff22110fdf32100fdf;
assign testcases[406] = 512'h50551dce60631cde52100fff51000fff40100fff40100dff40100fdf40100fdf62663bde52553cce32110fef33110eef44210dff43310dff22110fdf32100fdf;
assign testcases[407] = 512'h20100fef20100fff41000fff40000fff20000fff30000fff30000fef30000fef21110fff21110fef21000fff21000fff21000fff21000fff11000fef21000fef;
assign testcases[408] = 512'h20110fef30210eef41000fff50000fff20000fff30000fff30000fef30000fef21221eef21221eee21000fff21000fff22100fff22100fff21000fef21000fef;
assign testcases[409] = 512'h20220ede30210eef41000fff50000fff30000fff30000fff30000fef30000fef31321def31221ede21000fff21000fff22100fff32100fff21000fef21000fef;
assign testcases[410] = 512'h30221ede40320def41000fff50000fff30000fff30000fff30000fef40000fef41331dde31332dde21100fef21100fef32100fff32200eff21000fef21100fef;
assign testcases[411] = 512'h30331ede40320def41000fff50000fff30000fff30000fff40100fef40000fef41432cde41332dde21100fef31100fef32200eff32200eff21100fef21100fef;
assign testcases[412] = 512'h30331edf40420def51000fff50000fff30000fff40000eff40100fef40100fef41442cdf41442dde21100fef32100fef33200eff32200eff22100fef22100fef;
assign testcases[413] = 512'h40331dde50420cef52000fff50000fff30000fff40000eff40100fef40100fef52442cde42442dce31110fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[414] = 512'h40441dde50430cef52000fff50000fff30000fff40100eff40100fef40100fef52552cde42442dde31110fef32110fef33210eff33200eff22110fef22100fef;
assign testcases[415] = 512'h40441ddf50531cef52000fff50000fff30100fff40100eff40100fef40100fef52552cdf52553cde31110fef32110fef33210eff33200eff22110fef32100fef;
assign testcases[416] = 512'h40441dde50531cef52000fff50000fff30100fff40100eff40100fef40100fef52552bde52553cde31110fef32110fef33210eff43200eff22110fef32100fef;
assign testcases[417] = 512'h40441dde50531cdf52000fff50000fff30100fff40100eff40100fef40100fef62552bde52553cde31110fef32110fef43210eff43200eff22110fef32100fef;
assign testcases[418] = 512'h40451dce60531cde52000fff51000fff40100fff40100eff40100fef40100fef62663bce52553cce31110fef32110fef43210dff43310dff22110fef32100fef;
assign testcases[419] = 512'h50451dce60531bdf52000fff51000fff40100fff40100eff40100fef40100fef62663bce52553cce32110fef33110fef43210dff43210dff22110fef32100fdf;
assign testcases[420] = 512'h50551dde60641bef52100fff51000fff40100fff40100eff40100fef40100fef62663bdf52663cce32110fef32110fef43210dff43310dff22110fef32100fef;
assign testcases[421] = 512'h50551ddf60641bef52100fff51000fff40100fff40100dff40100fef40100fef62673bdf52663cce32110fef32110fef44310dff43310dff22110fef32100fef;
assign testcases[422] = 512'h10111fef20110fff41000fff40000fff20000fff20000fff30000fef30000fef20111fff10111fef20000fff21000fff21000fff21100fff10000fef21000fef;
assign testcases[423] = 512'h20110fef30210eef41000fff50000fff20000fff30000fff30000fef30000fef31211eef21211eee21000fff21000fff22100fff22100fff21000fef21000fef;
assign testcases[424] = 512'h20220ede30310eef41000fff50000fff20000fff30000fff30000fef30000fef31321def31221ede21000fff21000fff22100fff32100fff21000fef21000fef;
assign testcases[425] = 512'h30221ede40320def41000fff50000fff30000fff30000fff30000fef30000fef41331dde31332dde21000fff21100fef32100fff32200fff21000fef21100fef;
assign testcases[426] = 512'h30331edf40320def41000fff50000fff30000fff30000fff40100fef40000fef41442cde41332dde21100fef31100fef32200eff32200eff21100fef22100fef;
assign testcases[427] = 512'h30331edf40420def52000fff50000fff30000fff40000eff40100fef40100fef52442cdf42432ddf21100fef32100fef33200eff33200eff22100fef22100fef;
assign testcases[428] = 512'h40331dde50420cee51000fff50000fff30000fff40000eff40100fef40100fef51442cde41442dce21100fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[429] = 512'h40441dde50430cee52000fff50000fff30000fff40000eff40100fef40100fef51552cde41442dde31110fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[430] = 512'h40441dde50530cdf52000fff50000fff30000fff40000eff40100fef40100fef52552bde52442cde31110fef32110fef33200eff33200eff22110fef22100fef;
assign testcases[431] = 512'h40441dde50530cee52000fff50000fff30000fff40100eff40100fef40100fef62552bde52553cde31110fef32110fef33210eff43200eff22110fef22100fef;
assign testcases[432] = 512'h40441ddf60531cef52000fff51000fff30100fff40100eff40100fef40100fef62562bdf52553cde32110fef33110fef43210eff43310eff23110fef33100fef;
assign testcases[433] = 512'h40451dce60531cdf52000fff51000fff30100fff40100eff40100fef40100fef62663bde52553cce32110fef32110fef43210eff43310dff22110fef32100fef;
assign testcases[434] = 512'h50441dde60531cee52000fff51000fff40100fff40100eff40100fef40100fef62652bde52553cce32110fef32110fef43210dff43210dff22110fef32100fdf;
assign testcases[435] = 512'h50551dce60641bdf52100fff51000fff40100fff40100dff40100fef40100fef62663bdf52663cce32110fef32110fef44210dff43310dff22110fef32100fef;
assign testcases[436] = 512'h10110fef20110fff41000fff40000fff20000fff20000fff30000fef30000fef20110fff10111fef20000fff20000fff21000fff21100fff10000fef20000fef;
assign testcases[437] = 512'h30220ede30210def41000fff50000fff20000fff30000fff30000fef30000fef31321def31221ede21000fff21000fff22100fff22100fff21000fef21000fef;
assign testcases[438] = 512'h30221ede40320def41000fff50000fff30000fff30000fff30000fef30000fef41331def31332dde21000fff21100fff32100fff32200fff21000fef21100fef;
assign testcases[439] = 512'h20110fef20100fff41000fff40000fff20000fff30000fff30000fef30000fef21110fff21110fef20000fff21000fff21000fff21100fff11000fef21000fef;
assign testcases[440] = 512'h20110fef30210eef41000fff50000fff20000fff30000fff30000fef30000fef31221eef21221eef21000fff21000fff22100fff22100fff21000fef21000fef;
assign testcases[441] = 512'h30220edf30310def41000fff50000fff30000fff30000fff30000fef30000fef31321def31321ede21000fff21000fff22100fff32100fff21000fef21000fef;
assign testcases[442] = 512'h30221ede40320def41000fff50000fff30000fff30000fff30000fef30000fef41331ddf31332dde21100fff21100fef32100fff32200eff21000fef21100fef;
assign testcases[443] = 512'h30331edf40320def41000fff50000fff30000fff30000fff40100fef40000fef41442cde41332dde21100fef32100fef32200eff32200eff21100fef22100fef;
assign testcases[444] = 512'h40341dde50430cef51000fff50000fff30000fff40000eff40100fef40100fef52452cdf42452dde21110fef32110fef33200eff33200eff22100fef22100fef;
assign testcases[445] = 512'h10000fef10000fff41000fff50000fff30000fff30000fff30000fef30000fef10000fff10100fff21100fef21100fff32100fff32100fff21000fef21100fef;
assign testcases[446] = 512'h10110fef20110fff51000fff50000fff30100fff40100eff40100fef40100fef11110fff21111fef31110fef31110fef33210eff33310eff21110fef21100fef;
assign testcases[447] = 512'h20110eef20210eef52100fff50000fff40100fff50100dff40100fef40100fef21211eef21221ede31110fef32110fef43310dff43310dff22110fef22101fef;
assign testcases[448] = 512'h20220edf20210eef52100fff51000fff40100fff50100dff40110fef40110fef21221eef21321edf32211fef32110fef44310dff44410dff32110fef32201fef;
assign testcases[449] = 512'h20220edf30210eef52100fff61000fff50100fff60100dff40110fef40110fef21221eef31221ddf32211fef32210fef54410dff54410cff32210fef32201fdf;
assign testcases[450] = 512'h30221edf30320def63100eff61000fff50110fff60110cff50210edf50211edf31331def32332ddf42221eef43221eef65410cff65520bff33221edf33211edf;
assign testcases[451] = 512'h30331ddf30320def63100eff61000fff60110fff70110bff50211edf50211edf32432cdf42442cce43221eef43221edf66520bff65620aef43221edf43311edf;
assign testcases[452] = 512'h30331dcf40420cef63100def71000fff70110eff80110aff60211ddf60211ddf42442cdf42453cce43321edf44331ddf76520aff76620aef44321edf44311ecf;
assign testcases[453] = 512'h40441ccf40430cef74100def71000fff70110eff80210aef60311ddf60211ddf42442bdf52553bce53331ddf54331ddf77620aef877209ef44331dcf54312dcf;
assign testcases[454] = 512'h40441cce40530cdf74200cef71000eff80210eff902109ef70311ccf60311dcf52552bcf53563bbe54431ddf54331ddf886209ef877208ef55431dcf55412dcf;
assign testcases[455] = 512'h40451cce50531bdf74200cef81000eff80210effa02108ef70311ccf70311ccf52552bcf53663abe54431ccf55431ccf987208ef977208ef55431ccf55412ccf;
assign testcases[456] = 512'h50551cce50531bdf85200bef81100eff90210effa02108ef70411ccf70311ccf52663acf63664abe64431ccf65431ccf997318ef988207ef55431cbf65512cbf;
assign testcases[457] = 512'h50561bce50641bdf85200bef81100eff90210effb02107ef80421bbf70411bbf52673acf6379dabe64541ccf65431ccfa98317efa88307ef66541cbf66512cbf;
assign testcases[458] = 512'h50661bbe50641bdf85200bef81100effa0210dffb02106ef80421bbf80411bbf63673acf637749be65541bcf66531bcfaa8317efa98206ef66541bbf66512bbf;
assign testcases[459] = 512'h10000fef10000fff41000fff50000fff30000fff30000fff30100fef30100fef10000fff10100fff21100fff21100fff32200fff32200fff21110fef21100fef;
assign testcases[460] = 512'h10110fef20100fff51000fff50000fff30100fff40100eff40100fef40100fef11110fff21111fef31110fef31110fef33210eff33310eff21110fef21100fef;
assign testcases[461] = 512'h20110fef20110fff52100fff50000fff40100fff50100eff40100fef40100fef21111eef21211eef31110fef32110fef43310dff43310dff22110fef32101fef;
assign testcases[462] = 512'h20110edf20210eef52100fff61000fff40100fff50100dff40110fef40110fef21221eef21221ede32211fef32110fef44310dff54410dff32210fdf32201fdf;
assign testcases[463] = 512'h20220edf30210eef52100eff61000fff50100fff60100dff50210fef50110fef21221eef32321ddf32221fef32210fef54410dff54410cff32220fdf32201fdf;
assign testcases[464] = 512'h30221ede30320def63100eff61000fff60110fff70110cff50210edf50211edf32331def32332dde42221edf43221eef65510cff65510bff33221edf43211edf;
assign testcases[465] = 512'h30331ddf40320def63100dff61000fff60110fff70110bff60211edf50211edf42432cdf42442cce43321edf43321edf66520bff75620aff43321edf43311edf;
assign testcases[466] = 512'h30331dcf40420cef73100def71000fff70110eff80110aff60311ddf60211ddf42442cdf42443bce53331ddf54321ddf76620aef76620aef44331ddf44311dcf;
assign testcases[467] = 512'h40441ccf40430cef74200def71000fff70210eff902109ef60311ddf60311dcf42452bdf53553bce53331ddf54331ddf876209ef877209ef54331dcf54412dcf;
assign testcases[468] = 512'h40441ccf40530cdf74200cef71000eff80210eff902109ef70311ccf70311ccf52552bdf53563bbe54431ddf54431ddf887209ef877208ef55431dcf55412dcf;
assign testcases[469] = 512'h40451cce50531bdf84200cef81100eff80210effa02108ef70411ccf70311ccf52552bcf53663abe64431ccf65431cdf987218ef977208ef55431ccf55512ccf;
assign testcases[470] = 512'h50551cce50531bdf85200bef81100eff90210effa02107ef70421ccf70411ccf53663acf63664abe64441ccf65431ccf997318ef988207ef65541cbf65512cbf;
assign testcases[471] = 512'h50551bce50641bdf85210bef81100eff90210effb02107ef80421bbf80411bbf63663acf63774abe65542bcf66531bcfa98317efa88306ef66541bbf66512bbf;
assign testcases[472] = 512'h50561bbe50641bdf85210aef92100effa0210dffb02106ef80421bbf80411bbf63673acf637749be75542bcf66531bcfaa8317efa98306ef66541bbf66612bbf;
assign testcases[473] = 512'h10000fef10000fff41000fff50000fff30000fff30000fff30000fef40000fef10000fff10100fff21100fff21100fff32100fff32100fff21100fef21100fef;
assign testcases[474] = 512'h10110fef20100fff51000fff50000fff30100fff40100eff40100fef40100fef11110fff21111fef31110fef31110fef33210eff43210eff21110fef22100fef;
assign testcases[475] = 512'h20110fef20110fff52100fff50000fff40100fff50100dff40100fef40100fef21111eef21211eef31110fef32110fef43310dff43310dff22110fef32101fef;
assign testcases[476] = 512'h20110eef20210eef52100fff61000fff40100fff50100dff40110fef40110fef21221eef22221edf32211fef32210fef44310dff54410dff32210fef32201fef;
assign testcases[477] = 512'h20220edf30210eef52100eff61000fff50100fff60100dff50210eef50110fef21221eef32321ddf32221fef32220eef54410dff54410cff32220fdf32201fdf;
assign testcases[478] = 512'h30221edf30320def63100eff61000fff60110fff70110cff50210edf50211edf32331def32332ddf42221eef43221eef65510cff65510bff33221edf43311edf;
assign testcases[479] = 512'h30331ddf40320def63100def71000fff60110fff70110bff60211ddf60211edf42432cdf43442cce43321edf43321edf66520bef76620aff44321edf44311edf;
assign testcases[480] = 512'h40331dcf40420cef74100def71000fff70110eff80210aff60311ddf60211ddf42442cdf43553cce53331ddf54331ddf77620aef76620aef44331dcf44311dcf;
assign testcases[481] = 512'h40441ccf40430cef74200cef71000fff70210eff902109ef60311dcf60311dcf42552bdf53553bce53431ddf54331ddf876209ef877209ef55431dcf54412dcf;
assign testcases[482] = 512'h40441ccf50530bdf74200cef81100eff80210eff902109ef70311ccf70311ccf53552bdf53663bbe54431ddf55431cdf887209ef877208ef55431dcf55412dcf;
assign testcases[483] = 512'h40551cce50531bdf85200cef81100eff90210effa02108ef70411ccf70311ccf53552bcf64663abe64441ccf65431ccf987318ef988208ef55441ccf65512cbf;
assign testcases[484] = 512'h50551bce50531bdf85210bef81100eff90210effa02107ef70421bcf70411ccf53663acf64674abe64541ccf65431ccf997318ef988207ef66541cbf65512cbf;
assign testcases[485] = 512'h50551bce50641bdf85210bef81100eff90210effb02107ef80421bbf80421bbf63663acf64774abe65542bcf66541bcfa98317efa88206ef66541bbf66512bbf;
assign testcases[486] = 512'h50561bbe60641adf96210aef92100effa0210dffb02106ef80521bbf80421bbf63673acf647749ae75542bcf76541bcfaa8316efa99306ef66541bbf76612bbf;
assign testcases[487] = 512'h10000fef10000fff41000fff50000fff20000fff30000fff30100fef30000fef11000fff11100fff20100fff21100fff21100fff21200fff21100fef21100fef;
assign testcases[488] = 512'h10110fef20100fff51000fff50000fff30100fff40100eff40100fef40100fef11110fff21111fef31110fef31110fef33210eff43210eff22110fef22100fef;
assign testcases[489] = 512'h20110fef20110fff52100fff50000fff40100fff50100dff40100fef40100fef21111eef21221eef31110fef32110fef43310dff43310dff32110fef32101fef;
assign testcases[490] = 512'h20110eef20210eef52100fff61000fff40100fff50100dff40110fef40110fef21221eef22221edf32211fef32210fef44310dff54410dff32210fef32201fdf;
assign testcases[491] = 512'h20220edf30210eef52100eff61000fff50100fff60100dff50210edf50110fef22221eef32321ddf32221fef32220fef55410dff54410cff33220fdf32201fdf;
assign testcases[492] = 512'h30221edf30320def63100eff61000fff60110fff70110cff50210edf50211edf32331def32332ddf42221eef43221eef65510cff65510bff33221edf43311edf;
assign testcases[493] = 512'h30331ddf40320def63100def71000fff60110fff70110bff60211ddf60211edf42432cdf43442cce43321edf43321edf66520bff75620aff44321edf43311edf;
assign testcases[494] = 512'h40331dcf40420cef74100def71000fff70110eff80110aff60311ddf60211ddf42442cdf43553cce53331ddf54331ddf77620aef766209ef44331dcf44311dcf;
assign testcases[495] = 512'h40441ccf40430cef74200cef71000fff70210eff902109ef60311dcf60311dcf43552bdf53553bce53431ddf54331ddf876209ef877209ef55431dcf54412dcf;
assign testcases[496] = 512'h40441ccf50530cdf74200cef81100eff80210eff902109ef70311ccf70311ccf53552bdf53663bbe54431cdf55431cdf887209ef877208ef55431dcf55412ccf;
assign testcases[497] = 512'h40551cce50531bdf85200cef81100eff90210effa02108ef70421ccf70311ccf53562bcf64664abe64441ccf65431ccf987318ef988208ef55441ccf65512ccf;
assign testcases[498] = 512'h50551cce50531bdf85210bef81100eff90210effa02107ef80421bcf70421bcf53663acf64674abe64542ccf65431ccf998317ef988207ef66541cbf65512cbf;
assign testcases[499] = 512'h50551bbe50641bdf85210bef81100eff90210effb02107ef80421bbf80421bbf63663acf64774abe65542bcf66541bcfa98317efa88206ef66541bbf66512bbf;
assign testcases[500] = 512'h50561bbe60641adf96210aef92100effa0210dffb02106ef80521bbf80421bbf63673acf647749ae75542bcf76541bcfaa8316efa99206ef67541bbf76612bbf;
assign testcases[501] = 512'h10000fef10000fff41000fff50000fff30000fff30000fff40100fef40000fef10000fff11100fff21100fff21100fff32100fff32200fff21100fef21100fef;
assign testcases[502] = 512'h10110fef20100fff51000fff50000fff40100fff40100eff40100fef40100fef11110fff21111fef31110fef31110fef33210eff43310eff22110fef22100fef;
assign testcases[503] = 512'h20110fef20110fff52100fff50000fff40100fff50100dff40100fef40100fef21111eef21211eef31110fef32110fef43310dff43310dff32110fef32201fef;
assign testcases[504] = 512'h20110eef20210eff52100fff61000fff40100fff50100dff40110fef40110fef21221eef22221edf32211fef32210fef44310dff54410dff32210fdf32201fdf;
assign testcases[505] = 512'h20220edf30210eef62100eff61000fff50100fff60100cff50210edf50110edf22221eef32321ddf32221fef42220eef54410cff54410cff33221fdf33201edf;
assign testcases[506] = 512'h30221edf30320def63100eef61000fff60110fff70110bff50210edf50211edf32331ddf33332dcf42221edf43221edf65520bff65510bff43221edf43311edf;
assign testcases[507] = 512'h30331ddf40320def63100def71000fff60110fff70110bff60211ddf60211ddf42432cdf43442cce43321edf43321edf76520bef76620aff44331edf44311edf;
assign testcases[508] = 512'h40331ddf40420cef74200def71000fff70110eff80210aff60311ddf60311ddf43442cdf43553cce53331ddf54331ddf77620aef766209ef44331dcf54411dcf;
assign testcases[509] = 512'h40441cce40430cdf74200cef71000eff80210eff902109ef70311ccf60311dcf43552bdf53553bce53431ddf54331ddf876209ef877209ef55431dcf54412dcf;
assign testcases[510] = 512'h40441cce50530cdf74200cef81100eff80210eff902109ef70411ccf70311ccf53552bdf54663bbe54431cdf55431cdf887209ef977208ef55431ccf55412ccf;
assign testcases[511] = 512'h40551cce50531bdf85200bef81100eff90210effa02108ef70421ccf70311ccf53552bcf64663abe64441ccf65431ccf987318ef988208ef65541ccf65512ccf;
assign testcases[512] = 512'h50551cce50531bdf85210bef81100eff90210effb02107ef80421bbf80421bcf53663acf64674abe64542ccf65441bcfa98317ef988306ef66541cbf65512cbf;
assign testcases[513] = 512'h50561bbe50631bdf85210bef91100effa0210dffb02107ef80421bbf80421bbf63663acf63774abe64542bcf66541bcfa98317efa89316ef66541bbf66612bbf;
assign testcases[514] = 512'h50661bbe50641ade95210aef91100effa0210dffc02106ef80521bbf80421bbf63673ace637849ad75542bcf76541bcfb98317efa99315ef76641bbf76612baf;
assign testcases[515] = 512'h10000fef10000fff86310bef82100eff50110fff60110bff60421ccf60421ccf10000fff00000fff65542ccf56541ccf55410cff55410bff46441dcf55412dcf;
assign testcases[516] = 512'h10000fef10000fff86310aef92100eff60110fff70110bff70421ccf70421ccf10000fff00000fff65652ccf67541bcf56410bff66510aff56541dcf56512dcf;
assign testcases[517] = 512'h10000fef10000fff97310adf92100dff60110eff70110aef70521ccf70421ccf10000fff10000fff66652bcf67651bcf66520bef66510aef57552ccf56512ccf;
assign testcases[518] = 512'h10000fef10100fff984109df92100dff70110eff80110aef80521bbf80522bbf10000fff10000fff76762bbf78651abf67520aef76620aef57652cbf67612cbf;
assign testcases[519] = 512'h10000fef10100fffa84108dfa2100dff70110eff802109ef80631bbf80522bbf10000fff10000fff77763abf78762abf77520aef776209ef68662cbf67623cbf;
assign testcases[520] = 512'h10000fef10100fffa84108dfa2110dff70210eff802109ef80631abf80532abf10000fff10000fff87873abf897629bf786209ef776208ef68662bbf68723bbf;
assign testcases[521] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff40100fef40100fef00000fff00000fff21100fef31100fef21100fff21100fff21100fef21100fef;
assign testcases[522] = 512'h00000fff10000fff52100fff51000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef32100fff32200eff22110fef22100fef;
assign testcases[523] = 512'h10000fff10000fff63100eff61000fff30100fff40100eff40210fef40110fef00000fff00000fff32211fef33210fef33200eff33200eff33210fdf32201fef;
assign testcases[524] = 512'h10000fef10000fff63100eff61000fff40100fff40100eff50210edf50210edf00000fff00000fff43221eef43220eef33210eff43210eff33221fdf33201fdf;
assign testcases[525] = 512'h10000fef10000fff63200def61000fff40100fff50100dff50210edf50211edf00000fff00000fff43321edf44321eef43210eff43310dff33221edf33311edf;
assign testcases[526] = 512'h10000fef10000fff74200cef71100fff50100fff50100dff60311ddf60311ddf00000fff00000fff54431ddf54431ddf44310dff44310cff44331edf44311edf;
assign testcases[527] = 512'h10000fef10000fff75210cef81100eff50100fff60100cff60422ddf60322dcf00000fff00000fff54543ddf55442ddf55410cff55410cff45442dcf45413dcf;
assign testcases[528] = 512'h10000fef10000fff86310bef82100eff50100fff60110bff70421ccf70421ccf10000fff00000fff65542ccf66541ccf55410cff55510bff45441dcf55512dcf;
assign testcases[529] = 512'h10000fef10000fff96310aef92100eff60110fff70110bff70421ccf70421ccf10000fff00000fff65652bcf66541bcf66410bff66510bff56551dcf56512dcf;
assign testcases[530] = 512'h10000fef10000fff97310adf92100dff60110eff70110aef70521ccf70521bcf10000fff10000fff76762bcf77651bcf67520bef66510aef57552ccf56512ccf;
assign testcases[531] = 512'h10000fef10000fffa74109dfa2100dff70110eff801109ef80521bbf80522bbf10000fff10000fff76762abf78751abf67520aef776209ef67662cbf67613cbf;
assign testcases[532] = 512'h10000fef10100fffa84108dfa2100dff70210eff802109ef80631bbf80532bbf10000fff10000fff77873abf78762abf77520aef776209ef67662cbf67623cbf;
assign testcases[533] = 512'h10000fef10100fffa84108dfa2110dff70210eff902109ef80631abf80632abf11000fff11000fff878739bf897629bf786209ef876208ef68762bbf67723bbf;
assign testcases[534] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff40100fef40100fef00000fff00000fff21100fef31100fef21100fff21100fff21100fef21100fef;
assign testcases[535] = 512'h00000fff10000fff52100fff51000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef32100fff32200eff22110fef22100fef;
assign testcases[536] = 512'h10000fff10000fff62100eff61000fff30100fff40100eff40210fef40110fef00000fff00000fff32211fef32210fef33200eff33200eff32210fdf32201fef;
assign testcases[537] = 512'h10000fef10000fff63100eff61000fff40100fff40100eff50210edf50210edf00000fff00000fff42221eef43220eef33210eff33310eff33221fdf33201fdf;
assign testcases[538] = 512'h10000fef10000fff63100def61000fff40100fff50100dff50210edf50211edf00000fff00000fff43321edf43321eef43210eff43310dff33221edf33311edf;
assign testcases[539] = 512'h10000fef10000fff74200def71100fff40100fff50100dff60311ddf60311ddf00000fff00000fff53431ddf54431ddf44310dff44410cff44331edf44311edf;
assign testcases[540] = 512'h10000fef10000fff75210cef81100eff50100fff60100cff60421ddf60311dcf00000fff00000fff54541ddf55431ddf55410cff54410cff45431dcf44412dcf;
assign testcases[541] = 512'h10000fef10000fff85310bef82100eff50100fff60110bff70421ccf60421ccf10000fff00000fff65542ccf66541ccf55410cff55510bff45441dcf55512dcf;
assign testcases[542] = 512'h10000fef10000fff96310aef92100eff60110fff70110bff70521ccf70421ccf10000fff00000fff65652bcf66541bcf66410bff65510aff56552dcf55512dcf;
assign testcases[543] = 512'h10000fef10000fff97310adf92100dff60110eff70110aef70521bcf70521bcf10000fff00000fff76762bcf77651bcf66520bef66510aef56552ccf56512ccf;
assign testcases[544] = 512'h10000fef10000fff974109dfa2100dff70110eff80110aef80521bbf80522bbf10000fff10000fff76762abf77651abf67520aef766209ef57662cbf66612cbf;
assign testcases[545] = 512'h10000fef10100fffa84108dfa2100dff70210eff802109ef80631bbf80532bbf10000fff11000fff76873abf78762abf77520aef776209ef67662cbf67623cbf;
assign testcases[546] = 512'h10000fef10100fffa84108dfa2110cff80210eff902108ef80631abf80632abf11000fff11000fff878739bf887629bf786209ef876208ef68762bbf67723bbf;
assign testcases[547] = 512'h10000fef10100fffb94107dfb2110cff80210eff902108ef90631abf90632abf11100fff11000fff879739af898629af886209ef887208ef68772bbf78723bbf;
assign testcases[548] = 512'h10000fef10100fffa84108dfb2110cff80210eff902108ef80631abf90632abf11000fff10000fff878739bf888629af886209ef887208ef68762bbf67723baf;
assign testcases[549] = 512'h10000fef10100fffa64108dfa2110cff70210eff902108ef80632abf80632abf11000fff11000fff858739bf868729bf766209ef767208ef66772bbf65723baf;
assign testcases[550] = 512'h10451fef10531fffb84107dfb2100cff80210eff902108ef80721abf90621abf10563fff10664fff869529af888519af878319ef869317ef76852bbf66812baf;
assign testcases[551] = 512'h10000fef10100fffb75107dfb2110cff80210eff902108ef80632abe90632abe10100fff10100fff869839af888729af876209ef877208ef76772bbe66724bae;
assign testcases[552] = 512'h10000fef10000fff63200def71000fff40100fff50100dff50210edf50211edf00000fff00000fff43321edf43321eef43310eff43310dff33321edf33311edf;
assign testcases[553] = 512'h10000fef10000fff63200def71000fff40100fff50100dff50210edf50211edf00000fff00000fff43321edf43321eef43210eff43310dff33321edf33311edf;
assign testcases[554] = 512'h10000fef10000fff62200def71000fff40100fff40100dff50311edf50211edf00000fff00000fff42321edf42321edf32311eff42310dff32322edf32312edf;
assign testcases[555] = 512'h10000fef10000fff63200def71000fff40100fff50100dff50211edf50211edf00000fff00000fff42321edf43321edf43210dff43310dff33321edf33311edf;
assign testcases[556] = 512'h10000fef10000fff63200def71000fff40100fff50100dff50311edf50211edf00000fff00000fff43321edf43321edf43210eff43310dff33321edf33311edf;
assign testcases[557] = 512'h10000fef10000fff63200def71000fff40100fff50100dff50311edf50211edf00000fff00000fff43331edf43321edf43310dff43310dff33321edf33311edf;
assign testcases[558] = 512'h10000fef10100fffb85107cfb2110cff80210eff902108ef90632aaf90632aae11100fff11000fff879839ad898729ae886209ef887208ef78783baf77723baf;
assign testcases[559] = 512'h10000fef10100fffb85107dfb2110cff80210eff902108ef90632abf90632abf10000fff11000fff879839af888729af886208ef887208ef77773bbf77723bbf;
assign testcases[560] = 512'h10000fef10100fffb95107dfb3110cff80210eff902108ef90632abf90632abf11000fff11000fff889839af898729af886209ef887208ef78772bbf78723bbf;
assign testcases[561] = 512'h10000fef10000fffb85107dfb2110cff80210eff902108ef90632abf90632abf10000fff10000fff879839af988729af886208ef887208ef78772bbf77723bbf;
assign testcases[562] = 512'h10000fef10000fffa84108dfa2110dff80210eff902109ef80631bbf80532bbf10000fff00000fff86873abf88762abf776209ef776209ef67672bbf67623cbf;
assign testcases[563] = 512'h10000fef10000fffa74108dfa2110dff70210eff902109ef80631bbf80532bbf10000fff00000fff86873abf88762abf775209ef776209ef67672bbf66623cbf;
assign testcases[564] = 512'h10792fef20961fffab4108dfa3100dff80210eff902108ef80621abf80521abf219a4fff11895fef8a8529bf8c7419bf897209ef888208ef7c751bbf6b712baf;
assign testcases[565] = 512'h10210fef10210fffa94108dfa3100dff80210eff902108ef80631abf80522abf11221fff11221fff888739bf8a7619bf886209ef877208ef69762bbf68723baf;
assign testcases[566] = 512'h10000fff10000fff51000fff50000fff20000fff30000fff40100fef40100fef00000fff00000fff21110fef21110fff21100fff21100fff21110fef21100fef;
assign testcases[567] = 512'h10000fff10000fff52100fff51000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef22210fff32210fff22110fef22101fef;
assign testcases[568] = 512'h10000fef10000fff53100fff61000fff30100fff40100eff40110fef40110fef10000fff10000fff32211fef33210fef33210eff32210eff33210fef33201fef;
assign testcases[569] = 512'h10000fef10000fff63100eff61000fff30100fff40100eff40210fef50210fdf10000fff10000fff43221eef33220eef33210eff33210eff33220fdf33201fdf;
assign testcases[570] = 512'h10000fef10000fff63100eff61000fff40100fff50100eff50210edf50211edf10000fff10000fff43321eef43221eef43210eff43310dff33221edf33211edf;
assign testcases[571] = 512'h10000fef10100fff74200def71000fff40100fff50100dff50311edf50311edf10100fff10000fff53431ddf44331ddf44310dff44310dff44331edf44311edf;
assign testcases[572] = 512'h10000fef10100fff75210cef71100eff50100fff60100cff60311ddf60311ddf10100fff10000fff54541ddf55431ddf55310cff54410cff45431dcf45412dcf;
assign testcases[573] = 512'h10000fef10000fff85210bef81100eff50110fff60110bff60421dcf60421dcf10000fff10000fff64542ccf56541ccf55410cff55410bff55441dcf55412dcf;
assign testcases[574] = 512'h10000fef10000fff86310bef82100eff60110fff70110bff70421ccf70421ccf10000fff10000fff65652ccf66541ccf65410bff65510bff56541dcf56512dcf;
assign testcases[575] = 512'h10000fef10000fff86310aef92100eff60110fff70110bff70421ccf70421ccf10000fff10000fff65652bcf67541bcf66410bff65510aef56552ccf56512ccf;
assign testcases[576] = 512'h10000fef10000fff97310adf92100dff60110eff70110aff70521ccf70421ccf10100fff10000fff66652bcf68651bcf66510bef66520aef57552ccf57512cbf;
assign testcases[577] = 512'h10000fef10100fff983109df92100dff70110eff80110aef70521bbf80521bbf10100fff10000fff77762bbf78651abf77520aef775209ef68652cbf67612cbf;
assign testcases[578] = 512'h10000fef10100fff984109dfa2100dff70110eff802109ef80521bbf80522bbf10100fff10000fff77762abf79751abf77520aef776209ef68662cbf68623cbf;
assign testcases[579] = 512'h10220fef10210fffa94108dfa2100dff70210eff802109ef80521bbf80522abf11221fff11221fff87862abf79751abf786209ef776208ef69662bbf68623bbf;
assign testcases[580] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff40100fef40100fef00000fff00000fff21110fef21110fef21100fff21100fff21110fef21100fef;
assign testcases[581] = 512'h00000fff10000fff52100fff51000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef32100fff32200fff22110fef22100fef;
assign testcases[582] = 512'h10000fff10000fff53100eff61000fff30100fff40100eff40110fef40110fef00000fff00000fff32211fef33210fef33210eff32210eff33210fef33201fef;
assign testcases[583] = 512'h10000fef10000fff63100eff61000fff30100fff40100eff50210edf50210edf00000fff00000fff43221eef43220eef33210eff33210eff33221fdf33201fdf;
assign testcases[584] = 512'h10000fef10000fff64100eff61000fff40100fff50100eff50210edf50211edf10000fff00000fff43321eef44321eef43210eff43310dff33221edf33211edf;
assign testcases[585] = 512'h10000fef10000fff64200def71100fff40100fff50100dff50311edf50311edf10000fff10000fff43431ddf44331ddf44310dff44310dff44331edf44311edf;
assign testcases[586] = 512'h10000fef10000fff75200cef71100eff50100fff60100cff60311ddf60311ddf10000fff10000fff54431ddf55431ddf55310dff54410cff45431edf45411edf;
assign testcases[587] = 512'h10000fef10000fff76210cef82100eff50100fff60100cff60421dcf60311dcf10000fff10000fff55542ccf56441cdf55410cff55410cff46441dcf45412dcf;
assign testcases[588] = 512'h10000fef10000fff86310bef82100eff60110fff60110bff60421ccf70421ccf10000fff10000fff65542ccf67541ccf56410cff65410bff56441dcf56412dcf;
assign testcases[589] = 512'h10000fef10000fff87310bef92100eff60110fff70110bff70421ccf70421ccf10000fff10000fff66652bcf67541bcf66410bff66510aef57551dcf56512dcf;
assign testcases[590] = 512'h10000fef10000fff98310adf92100dff60110eff70110aff70521ccf70421ccf10000fff10000fff76652bcf68651bcf67510bef66520aef57552ccf57512cbf;
assign testcases[591] = 512'h10000fef10000fff983109df92100dff70110eff80110aef70521bbf80521bbf10000fff10000fff77762abf79651abf77520aef775209ef68652cbf68612cbf;
assign testcases[592] = 512'h10000fef10000fff994109dfa2100dff70110eff802109ef80521bbf80522bbf10000fff10000fff77762abf79761abf77520aef776209ef68662bbf68623bbf;
assign testcases[593] = 512'h10220fef10210fffa94108dfa3100dff80210eff902109ef80631abf80522abf11221fff11221fff888639bf8a7629bf786209ef877208ef69662bbf68723bbf;
assign testcases[594] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff40100fef40100fef00000fff00000fff21110fef31110fef21100fff21100fff21110fef21100fef;
assign testcases[595] = 512'h00000fff10000fff52100fff51000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef32100fff32200fff22110fef22100fef;
assign testcases[596] = 512'h10000fff10000fff53100eff61000fff30100fff40100eff40110fef40110fef00000fff00000fff32211fef33210fef33210eff32210eff33210fef33201fef;
assign testcases[597] = 512'h10000fff10000fff63100eff61000fff30100fff40100eff50210edf50210edf00000fff00000fff43221eef43220eef33210eff33210eff33221fdf33201fdf;
assign testcases[598] = 512'h10000fef10000fff63100eff61000fff40100fff40100eff50210edf50211edf00000fff00000fff43321eef43321eef33210eff43310dff33221edf33211edf;
assign testcases[599] = 512'h10000fef10000fff64200def71000fff40100fff50100dff50311edf50211edf10000fff00000fff43431ddf44331ddf44310dff44310dff44331edf44311edf;
assign testcases[600] = 512'h10000fef10000fff75210cef71100eff50100fff60100cff60311ddf60311ddf10000fff00000fff54431ddf55431ddf54310dff54410cff45431edf44411edf;
assign testcases[601] = 512'h10000fef10000fff75210cef81100eff50100fff60100cff60421dcf60321dcf10000fff00000fff54542ccf56441cdf55410cff55410cff45441dcf45412dcf;
assign testcases[602] = 512'h10000fef10000fff86310bef82100eff60110fff70110bff60421ccf70421ccf10000fff10000fff65542ccf66541ccf55410cff65410bff56441dcf56512dcf;
assign testcases[603] = 512'h10000fef10000fff86310bef82100eff60110fff70110bff70421ccf70421ccf10000fff10000fff65652bcf67541bcf66410bff66510aef56551dcf56512dcf;
assign testcases[604] = 512'h10000fef10000fff97310adf92100dff60110eff70110aff70521ccf70421ccf10000fff10000fff66652bcf67651bcf66510bef66520aef57552cbf56512cbf;
assign testcases[605] = 512'h10000fef10000fff973109df92100dff70110eff80110aef70521bbf80521bbf10000fff10000fff76762bbf78651abf77520aef765209ef67652cbf67612cbf;
assign testcases[606] = 512'h10000fef10000fff984109dfa2100dff70110eff802109ef80521bbf80522bbf10000fff10000fff77762abf79751abf77520aef776209ef68662cbf68623cbf;
assign testcases[607] = 512'h10210fef10210fffa94108dfa2100dff70210eff902109ef80621bbf80522abf11221fff11221fff87862abf897629bf786209ef776208ef68662bbf68623bbf;
assign testcases[608] = 512'h10441fef10530fff9c4109df93100dff70210eff802109ef80521bbf80521bbf11552fff11442fff7a762abf7d751abf79720aef787209ef6c662bbf6c723bbf;
assign testcases[609] = 512'h10110fef10110fff9a3109df93100dff70110eff801109ef80521bbf80521bbf11111fff10111fff79752abf7b651abf79510aef786109ef6a652bbf6a612bbf;
assign testcases[610] = 512'h00000fff10000fff41000fff50000fff20000fff30000fff30100fef30100fef00000fff00000fff21100fff21110fff21100fff21100fff21110fef21100fef;
assign testcases[611] = 512'h00000fff10000fff52000fff51000fff20000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef22100fff22100fff22110fef22100fef;
assign testcases[612] = 512'h10000fff10000fff53100fff51000fff30000fff40000fff40100fef40100fef00000fff00000fff32110fef33110fef33100fff33200eff23110fef23101fef;
assign testcases[613] = 512'h10000fef10000fff53100eff61000fff30100fff40100eff40110fef40110fef00000fff00000fff33211fef33210fef33210eff33210eff33210fef33201fef;
assign testcases[614] = 512'h10000fef10000fff53100eff61000fff30100fff40100eff40210fdf50210fdf00000fff00000fff33221eef34220eef33210eff33210eff34210fdf33201fdf;
assign testcases[615] = 512'h10000fef10000fff64100eff61000fff40100fff50100dff50210edf50211edf10000fff00000fff44321edf45321edf44210eff44310dff34221edf34311edf;
assign testcases[616] = 512'h10000fef10000fff65200def71000fff40100fff50100dff50311edf50211edf10000fff10000fff44431ddf45331ddf45310dff44310dff45331edf45311edf;
assign testcases[617] = 512'h10000fef10000fff76200cef72100eff50100fff60100cff60311ddf60311ddf10000fff10000fff55431ddf56431ddf55310dff55410cff46331edf46411ecf;
assign testcases[618] = 512'h10000fef10000fff77210cef82100eff50100fff60100cff60311dcf60311dcf10000fff10000fff56541ccf57431ccf56410cff56410bff47431dcf47412dcf;
assign testcases[619] = 512'h10000fef10000fff88310bef82100eff60110fff70110bff70421ccf70421ccf10000fff10000fff66542ccf68541ccf66410bff66510bff57441dcf57512dcf;
assign testcases[620] = 512'h10000fef10000fff88310adf92100dff60110eff70110aff70521ccf70421ccf10000fff10000fff66652bcf68651bcf67510bef66510aef57552ccf57512cbf;
assign testcases[621] = 512'h10000fef10000fff983109df92100dff70110eff80110aef70521bbf80521bbf10000fff10000fff77762abf79651abf77520aef776209ef68652cbf68612cbf;
assign testcases[622] = 512'h10000fef10000fffa94109dfa2100dff70210eff802109ef80531bbf80522bbf10000fff10000fff77762abf79762abf78520aef776209ef69662bbf68623bbf;
assign testcases[623] = 512'h10110fef10210fffaa4108dfa3100dff80210eff902109ef80621abf80522abf11221fff10211fff888629bf8a7629bf886209ef886208ef69662bbf69723bbf;
assign testcases[624] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff21100fff21110fef21100fef;
assign testcases[625] = 512'h00000fff10000fff52100fff51000fff30000fff40000fff40100fef40100fef00000fff00000fff32210fef32110fef32200fff32200fff22110fef22100fef;
assign testcases[626] = 512'h10000fff10000fff53100eff61000fff30100fff40100eff40210fef50110fef00000fff00000fff32211fef33210fef33210eff32210eff33210fef33201fef;
assign testcases[627] = 512'h10000fff10000fff63100eff61000fff40100fff40100eff50210edf50210edf00000fff00000fff43321eef43220eef33210eff33310eff33221fdf33201fdf;
assign testcases[628] = 512'h10000fff10000fff63100eff61000fff40100fff50100eff50210edf50211edf00000fff00000fff43321eef44321eef43210eff43310dff33221edf33311edf;
assign testcases[629] = 512'h10000fef10000fff74200def71100fff40100fff50100dff50311edf50311edf00000fff00000fff43431ddf44331ddf44310dff44310dff44331edf44311edf;
assign testcases[630] = 512'h10000fef10000fff75210cef71100eff50100fff60100cff60311ddf60311ddf10000fff00000fff54431ddf55431ddf54310dff54410cff45431edf45411edf;
assign testcases[631] = 512'h10000fef10000fff76210cef82100eff50100fff60100cff60321dcf60311dcf10000fff00000fff55541cdf56441cdf55410cff55410cff46441dcf45412dcf;
assign testcases[632] = 512'h10000fef10000fff86310bef82100eff50110fff60110bff60421ccf60421ccf10000fff00000fff65542ccf67541ccf56410cff55410bff56441dcf56512dcf;
assign testcases[633] = 512'h10000fef10000fff87310bef82100eff60110fff70110bff70421ccf70421ccf10000fff00000fff66652bcf67541bcf66410bff66510bff57541dcf57512dcf;
assign testcases[634] = 512'h10000fef10000fff97310adf92100dff60110eff70110aff70521ccf70421ccf10000fff10000fff76652bcf68651bcf67520bef66520aef57552ccf57512cbf;
assign testcases[635] = 512'h10000fef10000fff98310adf92100dff70110eff80110aef70521bbf70521bbf10000fff10000fff77762bbf78651bbf67520aef77520aef68652cbf57612cbf;
assign testcases[636] = 512'h10000fef10000fff993109df92100dff70110eff80110aef70521bbf80521bbf10000fff10000fff77762abf79651abf77520aef775209ef68652cbf68613cbf;
assign testcases[637] = 512'h10110fef10210fff993109df93100dff70110eff802109ef80521bbf80521bbf11221fff10221fff78762abf7a751abf78510aef786109ef69652bbf69612cbf;
assign testcases[638] = 512'h00000fff10000fff41000fff50000fff20000fff30000fff30100fef40000fef00000fff00000fff21100fff21100fff21100fff21100fff21100fef21100fef;
assign testcases[639] = 512'h00000fff10000fff52100fff51000fff30000fff30000fff40100fef40100fef00000fff00000fff32110fef32110fef22100fff22100fff22110fef22100fef;
assign testcases[640] = 512'h10000fff10000fff53100fff51000fff30000fff40000fff40100fef40100fef00000fff00000fff32210fef33110fef33100fff32200eff23110fef23100fef;
assign testcases[641] = 512'h10000fff10000fff53100eff61000fff30100fff40100eff40110fef40110fef00000fff00000fff33211fef33210fef33210eff33210eff33210fdf33201fdf;
assign testcases[642] = 512'h10000fef10000fff64100eff61000fff40100fff40100eff50210edf50210edf00000fff00000fff43221eef44220eef33210eff33210eff34221fdf33201fdf;
assign testcases[643] = 512'h10000fef10000fff64200def71000fff40100fff50100dff50210edf50211edf00000fff00000fff44321edf44321edf44310dff44310dff34321edf34311edf;
assign testcases[644] = 512'h10000fef10000fff75200def71100fff50100fff50100dff50311ddf60311ddf10000fff00000fff54431ddf55431ddf45310dff44310cff45331edf45311edf;
assign testcases[645] = 512'h10000fef10000fff76210cef72100eff50100fff60100cff60311dcf60311dcf10000fff00000fff55441ddf56431ddf55310cff55410cff46431dcf46412dcf;
assign testcases[646] = 512'h10000fef10000fff86210bef82100eff50110fff60110bff60421dcf60321dcf10000fff00000fff55542ccf57541ccf56410cff55410bff56441dcf56412dcf;
assign testcases[647] = 512'h10000fef10000fff87310bef82100eff60110fff70110bff70421ccf70421ccf10000fff00000fff66652ccf67541ccf66410bff66510bff57541dcf57512dcf;
assign testcases[648] = 512'h10000fef10000fff88310adf92100dff60110eff70110aff70421ccf70421ccf10000fff10000fff66652bcf68651bcf67410bef66510aef57551ccf57512cbf;
assign testcases[649] = 512'h10000fef10000fff98310adf92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77752bbf79651bbf77510aef77520aef68552cbf68612cbf;
assign testcases[650] = 512'h10000fef10000fff993109dfa2100dff70110eff801109ef80521bbf80522bbf10000fff10000fff77762abf79751abf77520aef776209ef68652cbf68623cbf;
assign testcases[651] = 512'h10110fef10210fffa94108dfa3100dff70210eff802109ef80521bbf80521bbf11221fff10211fff78762abf8a751abf786209ef786209ef69652bbf68613bbf;
assign testcases[652] = 512'h10110fef10110fff9a310adf93100dff60110eff80110aef70421bbf70421bbf11110fff10110fff78652bbf7b541bbf68520aef776209ef5a551cbf5a512cbf;
assign testcases[653] = 512'h10000fef10000fff993109df92100dff70110eff80110aef70521bbf70421bbf10100fff10000fff77652bbf79641abf78510aef775109ef69552cbf68512cbf;
assign testcases[654] = 512'h10000fef10000fff99310adf92100dff60110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf79651bbf67510aef775209ef58552cbf58512cbf;
assign testcases[655] = 512'h20100fef30100fff41000fff50000fff20000fff30000fff30000fef30000fef21110fff21100fff21000fff21000fff21000fff21000fff21000fef21000fef;
assign testcases[656] = 512'h30110fef30110eff41000fff50000fff30000fff30000fff30000fef30000fef31110fff31110fef21000fff21000fff21100fff21100fff21000fef21000fef;
assign testcases[657] = 512'h40110edf40110eef41000fff50000fff30000fff40000fff40000fef40000fef41111eef31111eef21000fff21000fff32100fff32100fff21000fef21000fef;
assign testcases[658] = 512'h40210ddf50210def51000fff50000fff30000fff40000fff40000fef40000fef51221def41211ddf31000fef31000fff32100fff32100fff21000fef21000fef;
assign testcases[659] = 512'h50221dde60310cef52000fff50000fff30000fff40000fff40000fef40000fef51221cdf51221dde31000fef32000fef32100fff32100eff21000fef21000fef;
assign testcases[660] = 512'h60321cce60310bdf52000fff50000fff40000fff50000eff40000fef40000fef61321cdf51321cce31100fef32100fef42100eff42100eff32100fef32100fef;
assign testcases[661] = 512'h60431cce70420bdf52000fff51000fff40000fff50000eff40100fef40100fef61431bdf61332cce32100fef32100fef43100eff43100eff32100fef32100fef;
assign testcases[662] = 512'h1029ffef10000fff40a00fff60241fff60210eff702107ef70748abf7074babf00000fff00000fff71aaf9af71a9f9af628318ef629317ef5189fbaf5182fbbf;
assign testcases[663] = 512'h00168fff10000fff40cefdaf40472ccf30210fff40210fff40632fef40632fef00000fff00000fff31983fef31872fef32620fff32720eff21772fef21723fef;
assign testcases[664] = 512'h10000fce10000fdf40a00fff75472eee80210eff902108df80632abf90632abf10000fff00000fff878839bf898729bf886209ef877208ef78772bbf78723bbf;
assign testcases[665] = 512'h10000fbb10000fcc91a0080f52241eef80210bb89021000080632a6090632a7410000fff00000fed8798395089872900876202008772000078772b8577723b52;
assign testcases[666] = 512'h1f110fef13210fffa2cf06cfcf583b73bf8efdffcf7cf7efafb7f9afafa6f9af10111fff10111fffa8cf88afaabd48afa9ffa7efa8efa6ef89af9aaf89ef8aaf;
assign testcases[667] = 512'h10000f9c10100d5cb37246cfc148400090431000a043174990a659af90a689af00110fff00000fff92bd88af93ab48af958417bf957206cf73772aaf73723aaf;
assign testcases[668] = 512'h00010fff00110fff41110fff40221fff20321fff30110fff30111fef30966fef00000fff00000fff41dd5edf41dd3edf52b31bef63b418ef529c5cbf52a48b9f;
assign testcases[669] = 512'h00000fff10100fff51720fff40000fff40421fff40321fff40b63fef50a64fef00110fff00000fff31fe6fef31ed4fef41d41eff31e41eff31df6fef31e48fef;
assign testcases[670] = 512'h00000fff00000fff40000fff40000fff10000fff20000fff30000fef30000fef00000fff00000fff20000fff20000fff10000fff10000fff10000fef10000fef;
assign testcases[671] = 512'h00000fff00000fff40000fff40000fff10000fff20000fff30000fef30000fef00000fff00000fff20000fff20000fff10000fff10000fff10000fef10000fef;
assign testcases[672] = 512'h00000fff00000fff40000fff40000fff10000fff20000fff30000fef30000fef00000fff00000fff20000fff20000fff10000fff10000fff10000fef10000fef;
assign testcases[673] = 512'h00000fff00000fff40000fff40000fff10000fff20000fff30000fef30000fef00000fff00000fff20000fff20000fff10000fff10000fff10000fef10000fef;
assign testcases[674] = 512'h00000fff00000fff40000fff40000fff10000fff20000fff30000fef30000fef00000fff00000fff20000fff20000fff10000fff10000fff10000fef10000fef;
assign testcases[675] = 512'h00000fff00000fff40000fff40000fff10000fff20000fff30000fef30000fef00000fff00000fff20000fff20000fff10000fff10000fff10000fef10000fef;
assign testcases[676] = 512'h00000fff00000fff40000fff40000fff10000fff20000fff30000fef30000fef00000fff00000fff20000fff20000fff10000fff10000fff10000fef10000fef;
assign testcases[677] = 512'h00000fff00000fff40000fff40000fff10000fff20000fff30000fef30000fef00000fff00000fff20000fff20000fff10000fff10000fff10000fef10000fef;
assign testcases[678] = 512'h10110fef10100fff41000fff50000fff30110fff30100fff30110fef40110fef11110fff11110fef21110fef21110fff32310eff32310eff21110fef21101fef;
assign testcases[679] = 512'h10110fef10100fff41000fff50000fff30100fff40100fff40100fef40100fef11110fff11110fff21110fef21110fef32310eff32310eff21110fef21101fef;
assign testcases[680] = 512'h20110fef20110fff52100fff50000fff40110fff40100eff40110fef40110fef21110fff21111fef31110fef32110fef43410eff43410dff22110fef32101fef;
assign testcases[681] = 512'h20110fef20210eff52100fff51000fff50110fff50100eff40110fef40110fef21221eef22221eef32211fef32210fef54410dff53410dff32210fef32201fef;
assign testcases[682] = 512'h20220edf20210eef52100fff61000fff50110fff50100dff40110fef40110fef22221eef32221edf32221fef32220fef54510cff54510cff32221fdf32201fdf;
assign testcases[683] = 512'h20220edf30210eef52100eff61000fff60110fff60110dff50210eef50111edf32221def32321ddf42221eef43220eef65520cff64520bff33221edf33211edf;
assign testcases[684] = 512'h30331ddf30320def63100eff61000fff70210eff70110cff50210edf50211edf32331ddf43332ddf43321edf43221edf75620bff75620aff44321edf43311edf;
assign testcases[685] = 512'h40331dcf40320cef63100dff61000fff70210eff70110bff50211edf60211edf43442cdf43442cce43331ddf54321ddf86720aef867209ef44331edf44311dcf;
assign testcases[686] = 512'h40441ccf40420cef64100def71000fff80210eff80110aff60311ddf60211ddf43542bdf53553bce53331ddf54331ddf877209ef868208ef55431dcf54411dcf;
assign testcases[687] = 512'h40441cce50430bdf74200def71000fff90210eff80210aef60311dcf60311dcf53552bdf53553bbe54431ddf55431cdf978208ef979308ef55431dcf55412dcf;
assign testcases[688] = 512'h50551bce50530bdf74200cef71000effa0210eff902109ef70311ccf70311ccf53562bcf63663abe64431ccf65431ccfa88318efa79317ef55431ccf65512cbf;
assign testcases[689] = 512'h50551bbe50531bdf75200cef81100effa0210dffa02108ef70311ccf70311ccf64663acf63664abe64531ccf66441ccfa89317efa8a316ef66541cbf66512cbf;
assign testcases[690] = 512'h50661bbe60631adf85200bef81100effb0210dffa02108ef70421ccf70311ccf64673acf64774abe65541bcf66541bcfb99317efb8a315ef66541bbf66512bbf;
assign testcases[691] = 512'h60662abe60641adf86210bef81100effb0310dffa02107ef70421bbf80411bcf647739cf747749ae75542bcf76541bcfb99316efb8a315ef77541bbf76612baf;
assign testcases[692] = 512'h10110fef10100fff41000fff50000fff30100fff40100fff40100fef40100fef11110fff11110fff21110fef21110fff32310eff32310eff21110fef21100fef;
assign testcases[693] = 512'h20110fef20110fff52100fff50000fff40100fff40100eff40100fef40100fef21110fff21111fef31110fef32110fef43310eff43410dff22110fef32101fef;
assign testcases[694] = 512'h20110fef20210eff52100fff51000fff50110fff50100eff40110fef40110fef21211eef21221eef32211fef32110fef54410dff53410dff32210fef32201fef;
assign testcases[695] = 512'h20220edf20210eef52100fff61000fff50110fff50100dff40110fef50110fef22221eef32221edf32211fef32210fef54410cff54510cff33210fdf33201fdf;
assign testcases[696] = 512'h30220edf30210eef52100eff61000fff60110fff60100dff50210edf50110edf32221def32321ddf42221eef43220eef65510cff64510bff33221edf33211edf;
assign testcases[697] = 512'h30331ddf30320def63100eff61000fff70210fff70110cff50210edf50211edf32331ddf42332cde43321eef43221eef75620bff75620aff44321edf44311edf;
assign testcases[698] = 512'h40331dcf40320cef63100eff71000fff80210eff70110bff60211edf60211edf43442cdf43442cce53321ddf54321ddf86720aef867209ef44321edf44311dcf;
assign testcases[699] = 512'h40441cce40420cef64100def71000fff80210eff80210aff60311ddf60211ddf43542bdf53553bce53331ddf54331ddf877209ef868208ef55431dcf55411dcf;
assign testcases[700] = 512'h40441cce50430bdf74200def71000fff90210eff90210aff60311dcf60311dcf53552bdf53553bbe54431ddf55431ddf978209ef979308ef55431dcf55412dcf;
assign testcases[701] = 512'h50551bce50530bdf74200cef71000effa0210eff902109ef70311ccf70311ccf53562bcf63663abe64431ccf65431ccfa88308efa79317ef55431ccf65512cbf;
assign testcases[702] = 512'h50551bbe50531bdf75200cef81100effa0210dffa02109ef70421ccf70311ccf64663acf64664abe64541ccf65441ccfa89317efa8a316ef66541cbf66512cbf;
assign testcases[703] = 512'h50661bbe60631adf85210bef81100effb0210dffa02108ef70421ccf70411ccf64673acf64774abe65541bcf66541bcfb99317efb8a315ef66541bbf66612bbf;
assign testcases[704] = 512'h60662abe60641adf85210bef81100effb0310dffb02107ef80421bbf80421bbf647739cf747749ae75542bcf76541bcfb99316efb8b315ef77641bbf76612bbf;
assign testcases[705] = 512'h10000fef10100fff41000fff50000fff30100fff40000fff40100fef40100fef11100fff11110fff21110fef21110fef32210eff32210eff21110fef21100fef;
assign testcases[706] = 512'h20110fef20110fff52000fff50000fff40100fff40100eff40100fef40100fef21110fff21111fef31110fef32110fef43310eff43310dff22110fef32100fef;
assign testcases[707] = 512'h20110fef20110eff52100fff51000fff50100fff50100dff40110fef40100fef22211eef22221eef32210fef32110fef54410dff53410cff32210fef32201fef;
assign testcases[708] = 512'h20220edf20210eef52100fff61000fff50110fff50100dff40110fef50110fef22221eef32221edf32211fef32210fef54410cff54510cff32210fdf32201fdf;
assign testcases[709] = 512'h30220edf30210eef52100eff61000fff60110fff60100dff50210edf50110edf32221def32321ddf42221eef43220eef65510cff64510bff33220edf33211edf;
assign testcases[710] = 512'h30331ddf30320def63100eff61000fff70210eff70110cff50210edf50211edf32331ddf42332cdf43321eef43221eef75620bff75720aff43321edf43311edf;
assign testcases[711] = 512'h40331dcf40320cef63100def71000fff80210eff70110bff60211ddf60211ddf43442cdf43442cce53331ddf54321ddf86720aef867209ef44331ddf44311dcf;
assign testcases[712] = 512'h40441ccf40420cef74100def71000fff80210eff80210aff60311ddf60311ddf43542bdf53553bce53431ddf54331ddf877209ef968208ef55431dcf54411dcf;
assign testcases[713] = 512'h40441cce50430bdf74200cef71000eff90210eff90210aff60311dcf60311dcf53552bdf54553bbe54431cdf55431cdf978308ef979308ef55431dcf55512ccf;
assign testcases[714] = 512'h50551bce50530bdf74200cef81100effa0210dff902109ef70311ccf70311ccf54662acf64663abe64441ccf65431ccfa88318efa79317ef65541ccf65512cbf;
assign testcases[715] = 512'h50551bbe50531bdf85200cef81100effa0210dffa02108ef70421ccf70311ccf64663acf64664abe64541ccf65441ccfa89317efa8a316ef66541cbf66512cbf;
assign testcases[716] = 512'h50561bbe60631adf85210bef81100effb0310dffa02108ef80421bcf80421bbf64673acf64774abe75542bcf76541bcfb99316efb8a315ef66541bbf76612bbf;
assign testcases[717] = 512'h60662bbe60641adf86210bef81100effb0310dffb02107ef80421bbf80421bbf647739cf747749ae75642bbf76541bbfb9a316efc8b315ef77641bbf76612baf;
assign testcases[718] = 512'h10100fef10100fff41000fff50000fff30100fff40100fff40100fef40100fef11110fff11110fff21110fef21110fef32310eff32310eff21110fef21100fef;
assign testcases[719] = 512'h20110fef20110fff52100fff50000fff40110fff40100eff40110fef40110fef21110fff21111fef31110fef32110fef43310dff43410dff22110fef32101fef;
assign testcases[720] = 512'h20110fef20110eff52100fff51000fff50110fff50100dff40110fef40110fef22211eef22221eef32211fef32210fef54410dff53510cff32210fef32201fdf;
assign testcases[721] = 512'h20220edf20210eef52100fff61000fff50110fff50100dff50210fef50110fef22221eef32221edf32221fef32220fef54510cff64510cff33221fdf33201fdf;
assign testcases[722] = 512'h20220edf30210eef52100eff61000fff60110fff60110cff50210edf50211edf32221def32321ddf42221eef43221eef65520cff64620bff33221edf33211edf;
assign testcases[723] = 512'h30331ddf30320def63100eff61000fff70210eff70110bff50211edf50211edf33331ddf43332ddf43321edf43321edf76620bff75720aff44321edf44311edf;
assign testcases[724] = 512'h40331dcf40320cef63100def71000fff80210eff80110bff60311ddf60211ddf43442cdf43442cce53331ddf54331ddf86720aef868209ef44331ddf54411dcf;
assign testcases[725] = 512'h40441ccf40420cef74200def71000fff90210eff80210aff60311dcf60311dcf43442bdf54553bce53431ddf54431ddf978209ef968208ef55431dcf55412dcf;
assign testcases[726] = 512'h40441cce50430bdf74200cef71000eff90210eff902109ef70311ccf70311ccf53552bdf54553bce64431ccf65431cdf978318ef979307ef55431ccf55512ccf;
assign testcases[727] = 512'h50551cce50530bdf74200cef81100effa0210dff902109ef70421ccf70311ccf54562bcf54663abe64541ccf65441ccfa89317efa7a316ef65541ccf65512cbf;
assign testcases[728] = 512'h50551bbe50531bdf85210bef81100effa0310dffa02108ef70421ccf70421ccf64663acf64664abe64542bcf65541bcfb89317efb8a316ef66541cbf66612bbf;
assign testcases[729] = 512'h50561bbe60631adf85210bef81100effb0310dffa02108ef80421bbf80421bbf64673acf64774abe75542bcf76541bcfb99316efb8a315ef66641bbf76612bbf;
assign testcases[730] = 512'h60661bbe60641adf85210aef91100effc0310dffb02107ef80421bbf80421bbf647739cf647749ae75642bbf76541abfc9a315efc8b314ef77651bbf76612baf;
assign testcases[731] = 512'h10000fef10100fff41000fff50000fff30100fff40100fff40100fef40100fef11100fff11110fff21110fef31110fef32210eff32310eff21110fef21100fef;
assign testcases[732] = 512'h20110fef20110fff51100fff50000fff40100fff40100eff40110fef40100fef21110fff21111fef31110fef32110fef43310dff43410dff22110fef32201fef;
assign testcases[733] = 512'h20110fef20110eff52100fff50000fff50110fff50100dff40110fef40110fef22211eef22221eef31211fef32210fef54410dff53410dff32210fef32201fef;
assign testcases[734] = 512'h20220edf20210eef52100fff61000fff50110fff50100dff40210fef50110fef22221eef32222edf32221fef32220fef54410cff54510cff32221fdf32201fdf;
assign testcases[735] = 512'h20220edf30210eef52100eff61000fff60110fff60110dff50210edf50211edf32221def32321ddf42221eef42220eef65520cff64520bff33221edf33211edf;
assign testcases[736] = 512'h30331ddf30320def63100eff61000fff70210fff60110cff50210edf50211edf32331ddf42332cde42321eef43221eef75620bff75620aff43321edf43311edf;
assign testcases[737] = 512'h40331dcf40320cef63100dff71000fff70210eff70110bff60211edf60211edf42442cdf42442cce43331ddf43321ddf76720aef867209ef44331edf44311dcf;
assign testcases[738] = 512'h40441ccf40420cef74100def71000fff80210eff80110aff60311ddf60211ddf42542bdf53553bce53331ddf54331ddf877209ef868209ef54431dcf54411dcf;
assign testcases[739] = 512'h40441cce50430bdf74200def71000fff90210eff80210aff60311dcf60311dcf52552bdf53553bbe54431ddf54431ddf978209ef978208ef55431dcf55412dcf;
assign testcases[740] = 512'h50551bce50530bdf74200cef81100effa0210eff902109ef70311ccf70311ccf53562acf63663abe64431ccf65431ccfa88308efa79307ef55431ccf65512cbf;
assign testcases[741] = 512'h50551bbe50531bdf85200cef81100effa0210dffa02108ef70421ccf70311ccf63663acf63664abe64541ccf65441ccfa89317efa79316ef65541cbf65512cbf;
assign testcases[742] = 512'h50561bbe60531adf85210bef81100effb0310dffa02108ef70421bcf70421bcf63673acf63774abe64542bcf65541bcfb89317efb8a316ef66541bbf66612bbf;
assign testcases[743] = 512'h60662abe60641adf85210bef81100effb0310dffb02107ef80421bbf80421bbf637739cf737749ae75542bcf76541bcfb99316efb8a315ef76641bbf76612bbf;
assign testcases[744] = 512'h10000fef10000fff98310adf92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf79651abf77510aef775109ef68552cbf68512cbf;
assign testcases[745] = 512'h10000fef10000fff993109df92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf79651abf78510aef775109ef58552cbf68512cbf;
assign testcases[746] = 512'h10000fef10000fff983109df92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf79651abf67510aef775109ef58552cbf68612cbf;
assign testcases[747] = 512'h10000fef10000fff993109df92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf79651abf67510aef775109ef58552cbf68512cbf;
assign testcases[748] = 512'h10000fef10000fff98310adf92100dff60110eff80110aef70521bbf70521bbf10000fff10000fff77652bbf78651abf67520aef775209ef58652cbf57612cbf;
assign testcases[749] = 512'h10000fef10000fff89310adf92100dff60110eff70110aef70421bbf70421bbf10000fff10000fff67652bcf69641bbf67410aef67510aef59551cbf58512cbf;
assign testcases[750] = 512'h10000fef10000fff99310adf92100dff70110eff80110aef70421bbf70421bbf10000fff10000fff77652bbf7a641abf78410aef775109ef69541cbf68512cbf;
assign testcases[751] = 512'h10000fef10000fff833109df91100dff60210eff70210aef70531bbf70522bbf10000fff10000fff63762bbf64662abf64520aef636209ef53662cbf53623cbf;
assign testcases[752] = 512'h10000fef10000fff983109df92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf78651abf77510aef775209ef58552cbf57612cbf;
assign testcases[753] = 512'h10000fef10000fff97310adf92100dff60110eff70110aef70521bbf70421bbf10000fff10000fff66652bbf77651abf67510aef665209ef56552cbf56512cbf;
assign testcases[754] = 512'h10000fef10000fff96310adf92100dff60110eff70110aef70521bbf70421bbf10000fff10000fff65652bbf66651bbf67510aef66510aef56551cbf55512cbf;
assign testcases[755] = 512'h10000fef10000fff99310adf92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf79651abf68510aef775109ef59552cbf58512cbf;
assign testcases[756] = 512'h10000fef10000fff993109df92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf79651abf78510aef775209ef68552cbf68612cbf;
assign testcases[757] = 512'h10000fef10000fff993109df92100dff70110eff80110aef70521bbf70421bbf10000fff10000fff77652bbf79651abf78510aef775209ef69552cbf68612cbf;
assign testcases[758] = 512'h10220fef10210fff9a4108dfa3100dff70210eff802109ef80621bbf80522bbf11321fff10221fff78862abf7a751abf786209ef787208ef69662bbf69723bbf;
assign testcases[759] = 512'h10110fef10110fff9a4109dfa3100dff70110eff802109ef80521bbf80521bbf11110fff10110fff78762abf7a751abf785209ef786209ef69652bbf69612bbf;
assign testcases[760] = 512'h10000fef10000fff8b310adf93100dff60110eff70110aef70421ccf70421cbf10000fff10000fff69652bcf6b641bcf68510aef68510aef5b541cbf5a512cbf;
assign testcases[761] = 512'h10000fef10000fff89310adf92100dff60110eff70110aef70421ccf70421bbf10000fff10000fff67642bbf69541bbf68410aef67510aef59541cbf58512cbf;
assign testcases[762] = 512'h10000fef10000fff86310adf92100dff60110eff70110aef70421bbf70421bbf10000fff00000fff65652bbf77651abf67510aef665109ef56552cbf56512cbf;
assign testcases[763] = 512'h10000fef10000fff98310adf92100dff70110eff80110aef70421bbf70421bbf10000fff00000fff77652bbf79651abf68510aef775109ef58551cbf68512cbf;
assign testcases[764] = 512'h10000fef10000fff993109df93100dff70110eff801109ef70521bbf80421bbf10000fff10000fff78652abf7a651abf78520aef775109ef69552cbf69612cbf;
assign testcases[765] = 512'h10000fef10000fff983109df92100dff70110eff801109ef80521bbf80521bbf10000fff00000fff77762abf78651abf77520aef776209ef68652bbf67612bbf;
assign testcases[766] = 512'h10100fef10100fffa94107dfb3110cff80210eff902108ef90631abf90632aaf11110fff10110fff889739af8a8629af886208ef887208ef79772baf79723baf;
assign testcases[767] = 512'h00000fff10000fff51000fff50000fff20000fff30000fff40100fef40100fef00000fff00000fff21110fef31110fef21100fff21100fff21110fef21100fef;
assign testcases[768] = 512'h00000fff10000fff52100fff61000fff30000fff40000fff40100fef40100fef00000fff00000fff32210fef32110fef32200fff32200eff22110fef32100fef;
assign testcases[769] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff50210fef50210fdf00000fff00000fff42221eef43220eef33210eff33210eff33210fdf33201fdf;
assign testcases[770] = 512'h10000fff10000fff63100eff61000fff40100fff50100dff50210edf50211edf00000fff00000fff43321eef43321eef43210eff43310dff33221edf33211edf;
assign testcases[771] = 512'h10000fff10000fff63200def71000fff40100fff50100dff50210edf50211edf00000fff00000fff43321edf44321edf43310dff43310dff33321edf43311edf;
assign testcases[772] = 512'h10000fef10000fff74210cef71100eff50100fff60100cff60311ddf60311ddf00000fff00000fff54441ddf54431ddf54410cff54410cff44431edf44411edf;
assign testcases[773] = 512'h10000fef10000fff85310bef81100eff60110fff70110bff60421dcf70421dcf00000fff00000fff64542ccf65541ccf55410cff64510bff55441dcf55512dcf;
assign testcases[774] = 512'h10000fef10000fff85310bef92100eff60110fff70110bff70421ccf70421ccf00000fff00000fff65652bcf66651bcf65520bff65520aef55552dcf55512dcf;
assign testcases[775] = 512'h10000fef10000fff96310adf92100dff70210eff80210aef70521ccf70522ccf10000fff00000fff75762bcf76651bcf76520aef75620aef66662ccf66613cbf;
assign testcases[776] = 512'h10000fef10000fff964109dfa2100dff70210eff802109ef80531bbf80522bbf10000fff00000fff75773abf77762abf76620aef766209ef66662cbf66623cbf;
assign testcases[777] = 512'h10000fef10000fffa74108dfa2110dff80210eff902109ef80631bbf80532abf10000fff00000fff86873abf88862abf876209ef867208ef67772bbf67723bbf;
assign testcases[778] = 512'h10000fef10000fffb84108dfb2110dff80210eff902108ef90632abf90632abf10000fff00000fff869839af888729bf876209ef877208ef77772bbf77723bbf;
assign testcases[779] = 512'h10000fef10000fffb85107dfb2110cff90210effa02107ef90732abf90632abf10000fff00000fff979839af989728af877208ef978207ef78883baf77824baf;
assign testcases[780] = 512'h00000fff10000fff51100fff50000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff32100fff21110fef21100fef;
assign testcases[781] = 512'h00000fff10000fff52100eff61000fff30100fff40100eff40110fef40110fef00000fff00000fff32211fef32210fef32210eff32210eff32210fef32201fef;
assign testcases[782] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff50210edf50211edf00000fff00000fff42321eef43221eef43210eff43310eff33221fdf33201fdf;
assign testcases[783] = 512'h10000fff10000fff63200dff71000fff40100fff50100dff50210edf50211edf00000fff00000fff43321edf43321eef43310dff43310dff33321edf33311edf;
assign testcases[784] = 512'h10000fff10000fff73200def71100fff50100fff50100dff50311edf60311edf00000fff00000fff53431ddf44331ddf43310dff43410dff43331edf43311edf;
assign testcases[785] = 512'h10000fef10000fff74210cef81100eff50100fff60110cff60321ddf60311ddf00000fff00000fff54541ddf54431ddf54410cff54410cff44441ddf44412dcf;
assign testcases[786] = 512'h10000fef10000fff85310bef81100eff60110fff70110bff70421ccf70421ccf00000fff00000fff64652ccf65541ccf65410cff64510bff55541dcf55512dcf;
assign testcases[787] = 512'h10000fef10000fff96310aef92100eff60110eff70110aff70521ccf70421ccf00000fff00000fff65652bcf66651bcf65520bef65520aef55552ccf55512ccf;
assign testcases[788] = 512'h10000fef10000fff96310adf92100dff70110eff80210aef70521bcf80522bcf10000fff00000fff75762bbf76651bcf76520aef75620aef66662cbf66623cbf;
assign testcases[789] = 512'h10000fef10000fffa74109dfa2100dff70210eff802109ef80531bbf80532bbf10000fff00000fff75873abf77762abf76620aef766209ef66662cbf66623cbf;
assign testcases[790] = 512'h10000fef10000fffa74108dfa2110dff80210eff902109ef80631bbf80632abf10000fff00000fff86873abf878729bf866209ef867208ef67772bbf66723bbf;
assign testcases[791] = 512'h10000fef10000fffb74108dfb2110cff80210eff902108ef90632abf90632abf10000fff00000fff869839af888729bf876209ef877208ef77772bbf77723bbf;
assign testcases[792] = 512'h10000fef10000fffb85107dfb2110cff90210effa02108ef90632aaf90632aaf10000fff00000fff979839af989728af877208ef977207ef78783baf77824baf;
assign testcases[793] = 512'h00000fff10000fff51100fff50000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff31200fff21110fef21100fef;
assign testcases[794] = 512'h00000fff10000fff52100eff61000fff30100fff40100eff40210fef40110fef00000fff00000fff32211fef32210fef32210eff32210eff32210fef32201fef;
assign testcases[795] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff50210edf50210edf00000fff00000fff42321eef43221eef33210eff43310eff33221fdf33201fdf;
assign testcases[796] = 512'h10000fff10000fff63200def71000fff40100fff50100dff50210edf50211edf00000fff00000fff43321edf43321edf43310dff43310dff33321edf33311edf;
assign testcases[797] = 512'h10000fff10000fff73200def71100fff40100fff50100dff50311edf50311edf00000fff00000fff43431ddf44331ddf43310dff43410dff43331edf43311edf;
assign testcases[798] = 512'h10000fef10000fff74210cef81100eff50110fff60110cff60321ddf60311ddf00000fff00000fff54541ddf54441ddf54410cff54410cff44441ddf44412ddf;
assign testcases[799] = 512'h10000fef10000fff85310bef81100eff60110fff70110bff60421dcf70421ccf00000fff00000fff64652ccf65541ccf55410cff64510bff55541dcf55512dcf;
assign testcases[800] = 512'h10000fef10000fff96310aef92100eff60110fff70110bff70521ccf70421ccf00000fff00000fff65652bcf66651bcf65520bff65520aff55552dcf55512dcf;
assign testcases[801] = 512'h10000fef10000fff96310adf92100dff70110eff80210aef70521bcf80522bcf10000fff00000fff75762bcf76651bcf76520aef75620aef66662ccf66623cbf;
assign testcases[802] = 512'h10000fef10000fffa74109dfa2100dff70210eff802109ef80531bbf80532bbf10000fff00000fff75873abf77762abf76620aef766209ef66662cbf66623cbf;
assign testcases[803] = 512'h10000fef10000fffa74108dfa2110dff80210eff902109ef80631bbf80532bbf10000fff00000fff86873abf87862abf876209ef867208ef67772bbf66723bbf;
assign testcases[804] = 512'h10000fef10000fffa74108dfb2110dff80210eff902108ef80632abf90632abf10000fff00000fff869839bf888729bf876209ef867208ef77772bbf77723bbf;
assign testcases[805] = 512'h10000fef10000fffb85107dfb2110cff80210effa02108ef90632aaf90632aaf10000fff00000fff979839af988729af877208ef977207ef77783baf77724baf;
assign testcases[806] = 512'h00000fff10000fff51100fff50000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff21100fff21110fef21100fef;
assign testcases[807] = 512'h00000fff10000fff52100fff61000fff30100fff40100eff40210fef40110fef00000fff00000fff32211fef32210fef32210eff32210eff32210fef32201fef;
assign testcases[808] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff50210edf50211edf00000fff00000fff42321eef43221eef33210eff42310eff32221fdf32201fdf;
assign testcases[809] = 512'h10000fff10000fff63200def71000fff40100fff50100dff50210edf50211edf00000fff00000fff42321edf43321edf43310dff43310dff33321edf33311edf;
assign testcases[810] = 512'h10000fff10100fff73200def71100fff40100fff50100dff50311edf50311edf00100fff00000fff53431ddf43331ddf43310dff43310dff43331edf43311edf;
assign testcases[811] = 512'h10000fef10000fff74210cef81100eff50110fff60110cff60321ddf60311dcf00000fff00000fff54541ddf54441ddf54410cff54410cff44441dcf44412dcf;
assign testcases[812] = 512'h00341fef10431fffc8fa16cfb2440cff90ff5dffb0ff66ef90ffa9afa0ffd9af11445fff10345fffa7ba48af99b928af989317ef97a316ef88993aaf78924aaf;
assign testcases[813] = 512'h10000fef10000fffb75107dfa2110dff90210effa02107ef90632abf90632abf10000fff00000fff969839af979828af877208ef968207ef76883baf76824baf;
assign testcases[814] = 512'h10000fef10000fffb85107dfa2110dff90210effa02107ef90732abf90632aaf10000fff00000fff969939af989828af877208ef978207ef77883baf77824baf;
assign testcases[815] = 512'h10000fef10000fffb85107cfb2110cff90210effa02107ef90732aae90632aaf10000fff00000fff969939ae989828af877208ef978207ef77883baf77824baf;
assign testcases[816] = 512'h10220fef10210fffc95106cfb2110cff90210dffb02106ef907429afa07429af11211fff11111fff97ba48af99a828af988217ef979206ef88993aaf78924aaf;
assign testcases[817] = 512'h10110e5f10110fffc65106cfb211035690210dffb02106ef907429afa07329af10110fff10000fff95a9489f97a827af977207ef978206ef76893aaf76824aaf;
assign testcases[818] = 512'h10000fef10000fffb75107df92110dff90210effa02107ef90732abf90632aaf10000fff00000fff969939af989828af977208ef978207ef77883baf77824baf;
assign testcases[819] = 512'h10000fef10000fffb75107cd92110dff90210effa02107ef90732aad90632aae10000fff00000fff9699399d9798289e877218ef978217ef76883bae76824bae;
assign testcases[820] = 512'h10000fef10000fffb85107dfa3110dff90210effa02107ef90732abf90632aaf10000fff00000fff969939af989828af977208ef978207ef77883baf77824baf;
assign testcases[821] = 512'h10000fef10000fffb85107dfa2110dff90210effa02107ef90732abf90632aaf10000fff00000fff969939af989828af977208ef978207ef77883baf77824baf;
assign testcases[822] = 512'h10110fef10210fffc85106cfa3110dff90210dffb02106efa07429afa07429af10211fff10111fffa7ba48afa9a827af988207efa79206ef88993aaf88924aaf;
assign testcases[823] = 512'h10110fef10110d7ec851064fa211068890210dffb02106ef907429afa07429af10110fff10100fffa7a9489fa9a827af988207efa79206ef88893aaf87824aaf;
assign testcases[824] = 512'h10000fff10000fff40bfffff52ffffff80210fff90210fff90632fef90633fef10000fff00000fff85984fff86973fff86720fff86720fff75783fef75724fef;
assign testcases[825] = 512'h00000fef10000fff40b00f6f40121fff6058aeff7047c8ef70423abf70424abf00000fff00000fff616549af616529af62eff8ef62eff7ef51562bbf51522baf;
assign testcases[826] = 512'h10000fef10000fff40000fff40000fff80210effa02108ef90632abf90632abf10000fff00000fff869839af989729af877208ef977207ef77783baf77724baf;
assign testcases[827] = 512'h10000fef10000fff40000fff40000fff80210effa02108ef90632abf90632abf10000fff00000fff979839af989729af877208ef978207ef78783bbf77724baf;
assign testcases[828] = 512'h10110fef10210fff40000fff63121fff90210dffb02107ef907429afa07329af10111fff10111fff97a948af99a828af987207ef988206ef88883aaf78824aaf;
assign testcases[829] = 512'h10110fef10100fff40000fff87110eff90210dffa02107ef907429afa07329af10110fff10000fff97a948af99a828af987207ef978206ef78883aaf78824aaf;
assign testcases[830] = 512'h10100fef10100fff40000fff87111eee90210dffb02107ef907429afa07329af10110fff10000fff97a938af999828af987207ef988206ef78883aaf78824aaf;
assign testcases[831] = 512'h10100fef10100fff40000a2f75111dce90210dffb02107ef907429afa07329af10110fff10000fff97a948af999828af987207ef978206ef78883aaf78824aaf;
assign testcases[832] = 512'h10000fef103fffff40a0081040342fde80210eff902108ef80631abf80632abf00000fff00000fff828739af838729af756208ef847208ef63772baf62723bbf;
assign testcases[833] = 512'h10231fef10320fff95310ade91100dff80210eff802109ef70521bbe70522bbf11331fff10221fff74873abe75762abf767209ef768208ef65772caf65723caf;
assign testcases[834] = 512'h10000fef10100fff973109df92100dff90210eff802109ef70521bbf80522bbf10100fff10000fff76873abf77762abf776209ef877208ef66662bbf66623cbf;
assign testcases[835] = 512'h10000fef10100fff983109df92100dff90210eff802109ef80521bbf80522bbf10100fff00000fff76873abf78762abf776209ef876208ef67662bbf67623cbf;
assign testcases[836] = 512'h10000fef10100fff983109df92100dff90210eff802109ef80521bbf80522bbf10000fff00000fff87873abf88762abf776209ef876208ef67662bbf67623cbf;
assign testcases[837] = 512'h10441fef10530fffa94108dfa2110dff90310dff902108ef80631abf80632abf10542fff10442fff879839af899729af888208ef889207ef78872baf78823baf;
assign testcases[838] = 512'h10110fef10110fffa74108dfa2100dff90210dff902108ef80631abf80522abf10110fff10110fff868739af888729af886208ef877207ef77772baf77723baf;
assign testcases[839] = 512'h10110fef10110fffa94108dfa2100dff90210dff902108ef80631abf80532abf10110fff10110fff878739af898729af886208ef887207ef78772baf78723baf;
assign testcases[840] = 512'h10110fef10100fffa94108dfa2100dff90210dff902108ef80631abf80532abf10110fff10110fff878739af898729af886208ef887207ef78772baf78723baf;
assign testcases[841] = 512'h10000fef10000fff953109dfa1100dff80210eff802109ef80521bbf80522bbf10000fff00000fff74862abf857629bf766209ef766208ef65662bbf65623bbf;
assign testcases[842] = 512'h10000fef10000fff984109dfa2100dff90210eff802109ef80521bbf80522bbf10000fff00000fff86873abf887629bf776209ef876208ef67662bbf67623bbf;
assign testcases[843] = 512'h10000fef10000fff984109dfa2100dff90210eff802109ef80521bbf80522bbf10000fff00000fff86873abf887629bf776209ef876208ef67662bbf67623bbf;
assign testcases[844] = 512'h10000fef10000fff984109dfa2100dff90210eff802109ef80531bbf80522bbf10000fff00000fff86873abf888629bf776209ef876208ef67662bbf67623bbf;
assign testcases[845] = 512'h10110fef10210fffa74108dfa2100dff90210dff902109ef80631abf80632abf11211fff11111fff869739af888729af876208ef877207ef77772baf76723baf;
assign testcases[846] = 512'h10100fef10100fffa64108dfa2100cff90210dff902108ef80631abf80532abf10110fff10000fff858739af868729af876208ef877207ef75772baf75723baf;
assign testcases[847] = 512'h10110fef10100fffa94108dfa2100cff90210dff902108ef80631abf90632aaf10110fff10100fff879739af898729af886208ef887207ef78772baf78723baf;
assign testcases[848] = 512'h10100fef10100fffa94108dfa2100cff90210dff902108ef80631abf90632abf10110fff10000fff879739af898729af886208ef887207ef78772baf78723baf;
assign testcases[849] = 512'h00000fff10000fff51000fff50000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff22100fff21110fef21100fef;
assign testcases[850] = 512'h00000fff10000fff52100fff51000fff30100fff30000fff40100fef40100fef00000fff00000fff32210fef32210fef32200fff32200eff22110fef22100fef;
assign testcases[851] = 512'h00000fff10000fff53100eff61000fff40100fff40100eff40210fef40110fef00000fff00000fff32221eef33220eef33210eff33210eff33210fdf33201fdf;
assign testcases[852] = 512'h10000fff10000fff63100eff61000fff40100fff40100eff50210edf50210edf00000fff00000fff43321eef43221eef33210eff43310eff33221fdf33211fdf;
assign testcases[853] = 512'h10000fff10000fff63100eff61000fff40100fff40100dff50210edf50211edf00000fff00000fff43321edf44321edf43310dff43310dff33321edf33311edf;
assign testcases[854] = 512'h10000fef10000fff74200def71100fff50110fff50100dff50311edf50311edf00000fff00000fff54431ddf55431ddf44310dff44410cff44331edf44311edf;
assign testcases[855] = 512'h10000fef10000fff75210cef71100eff60110fff60100cff60321dcf60311ddf00000fff00000fff54542ddf55441cdf55410cff54410cff45441dcf45412dcf;
assign testcases[856] = 512'h10000fef10000fff86210bef82100eff60110eff60110cff60421dcf60321dcf00000fff00000fff65552ccf66541ccf55410cff65510bff56441dcf56412dcf;
assign testcases[857] = 512'h10000fef10000fff86310bef82100eff70210eff70110bff70421ccf70421ccf10000fff00000fff65652bcf67651bcf66410bef66510aef56552dcf56512dcf;
assign testcases[858] = 512'h10000fef10000fff97310adf92100dff70210eff70110bff70521ccf70421ccf10000fff00000fff76762bcf77651bcf66520aef76620aef57552cbf57512ccf;
assign testcases[859] = 512'h10000fef10000fff97310adf92100dff80210eff70110aff70521ccf70522bbf10000fff00000fff76762abf78762abf77520aef766209ef67662cbf67623cbf;
assign testcases[860] = 512'h10000fef10000fff984109dfa2100dff80210eff80110aef80521bbf80522bbf10000fff00000fff77873abf78762abf77520aef776209ef68662cbf67623cbf;
assign testcases[861] = 512'h10000fef10000fffa84108dfa2100dff80210eff802109ef80531bbf80532bbf10000fff00000fff878739bf898629bf776209ef876208ef68772bbf68623bbf;
assign testcases[862] = 512'h00000fff10000fff52000fff50000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff22100fff21110fef21100fef;
assign testcases[863] = 512'h00000fff10000fff52100fff51000fff30100fff30000fff40100fef40100fef00000fff00000fff32210fef32210fef32200fff32200eff22110fef32101fef;
assign testcases[864] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff40210fef40110fef00000fff00000fff32221eef43220eef33210eff33210eff33220fdf33201fdf;
assign testcases[865] = 512'h10000fff10000fff63100eff61000fff40100fff40100eff50210edf50211edf00000fff00000fff43321eef43321eef33210eff43310dff33221fdf33211fdf;
assign testcases[866] = 512'h10000fff10000fff63100eff61000fff40100fff50100eff50210edf50211edf00000fff00000fff43321edf44321edf43310eff43310dff34321edf33311edf;
assign testcases[867] = 512'h10000fef10000fff75200def71100fff50110fff50100dff50311edf60311ddf00000fff00000fff54431ddf55431ddf44310dff54410cff44331edf44311edf;
assign testcases[868] = 512'h10000fef10000fff75210cef81100eff60110fff60100cff60321ddf60311ddf00000fff00000fff54542ddf55441cdf55410cff54410cff45441dcf45412dcf;
assign testcases[869] = 512'h10000fef10000fff86310bef82100eff60110eff60110cff60421dcf60421ccf00000fff00000fff65652ccf66541ccf55410cff65510bff56541dcf56512dcf;
assign testcases[870] = 512'h10000fef10000fff86310bef82100eff70210eff70110bff70421ccf70421ccf10000fff00000fff65652bcf67651bcf66410bef65510aff56552dcf56512dcf;
assign testcases[871] = 512'h10000fef10000fff97310adf92100dff70210eff70110bff70521ccf70421ccf10000fff00000fff76762bcf77651bcf66520bef66520aef57552ccf56512ccf;
assign testcases[872] = 512'h10000fef10000fff973109df92100dff80210eff70110aff70521bbf70522bbf10000fff00000fff76763abf78762abf77520aef766209ef67662cbf67623cbf;
assign testcases[873] = 512'h10000fef10000fff984109dfa2100dff80210eff80110aef80521bbf80522bbf10000fff00000fff77873abf78762abf77520aef776209ef68662cbf67623cbf;
assign testcases[874] = 512'h10000fef10000fffa84108dfa2100dff80210eff801109ef80531bbf80532bbf10000fff00000fff878739bf898629bf776209ef876208ef68672bbf68623bbf;
assign testcases[875] = 512'h00000fff10000fff51000fff50000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff22100fff21110fef21100fef;
assign testcases[876] = 512'h00000fff10000fff52100fff51000fff30100fff40000fff40110fef40100fef00000fff00000fff32210fef32210fef32200fff32200eff22110fef32101fef;
assign testcases[877] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff40210fef40110fef00000fff00000fff32221eef43220eef33210eff33210eff33220fdf33201fef;
assign testcases[878] = 512'h10000fff10000fff63100eff61000fff40100fff40100eff50210edf50211edf00000fff00000fff43321eef43321eef33210eff43310eff33221fdf33211fdf;
assign testcases[879] = 512'h10000fff10000fff63100def61000fff40100fff50100eff50210edf50211edf00000fff00000fff43321edf43321edf43310eff43310dff33321edf33311edf;
assign testcases[880] = 512'h10000fef10000fff74200def71100fff50110fff50100dff50311edf50311ddf00000fff00000fff53431ddf54431ddf44310dff54410cff44331edf44311edf;
assign testcases[881] = 512'h10000fef10000fff75210cef71100eff60110fff60100cff60311ddf60311dcf00000fff00000fff54542cdf55541cdf55410cff54410cff45441dcf44412dcf;
assign testcases[882] = 512'h10000fef10000fff85310bef81100eff60110eff60110cff60421dcf60421dcf00000fff00000fff64652ccf66541ccf55410cff65510bff55541dcf55512dcf;
assign testcases[883] = 512'h10000fef10000fff86310bef82100eff70210eff70110bff70421ccf70421ccf10000fff00000fff65652bcf66651bcf66410bff65510aff56552dcf56512dcf;
assign testcases[884] = 512'h10000fef10000fff87310adf92100dff70210eff70110bff70521ccf70421ccf10000fff00000fff76762bcf77651bcf66520bef66520aef57552ccf56512cbf;
assign testcases[885] = 512'h10000fef10000fff973109df92100dff80210eff70110aff70521bbf70522bbf10000fff00000fff76762abf78762abf76520aef766209ef67662cbf67623cbf;
assign testcases[886] = 512'h10000fef10000fff984109dfa2100dff80210eff80110aef80531bbe80522baf10000fff00000fff76873aaf88762aaf776209ef776209ef67662bbf67623bbf;
assign testcases[887] = 512'h10000fef10000fffa84108dfa2110dff80210eff802109ef80631bbf80532abf10000fff00000fff878739bf898629bf776209ef877208ef68772bbf68723bbf;
assign testcases[888] = 512'h00000fff10000fff51000fff50000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff21100fff21110fef21100fef;
assign testcases[889] = 512'h00000fff10000fff52100fff61000fff30100fff40000fff40110fef40110fef00000fff00000fff32211fef32210fef32210fff32210eff32210fef32201fef;
assign testcases[890] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff40210fef50210fdf00000fff00000fff42221eef43220eef33210eff33210eff33221fdf33201fdf;
assign testcases[891] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff50210edf50211edf00000fff00000fff43321eef43321eef43210eff43310dff33221edf33211edf;
assign testcases[892] = 512'h10000fff10000fff64200def61000fff40100fff50100dff50210edf50211edf00000fff00000fff43331edf44321edf43310dff43310dff34321edf33311edf;
assign testcases[893] = 512'h10000fef10000fff74200def71100fff50110fff50100dff60311ddf60311ddf00000fff00000fff54431ddf55431ddf44310dff54410cff44431edf44411edf;
assign testcases[894] = 512'h10000fef10000fff75210cef81100eff60110fff60100cff60321dcf60321dcf00000fff00000fff54542cdf55541cdf55410cff55410bff45441dcf45412dcf;
assign testcases[895] = 512'h10000fef10000fff86310bef82100eff60110eff60110cff60421ccf70421ccf00000fff00000fff65652ccf66541ccf65410bff65510bff56551dcf55512dcf;
assign testcases[896] = 512'h10000fef10000fff86310aef92100eff70210eff70110bff70421ccf70421ccf10000fff00000fff65652bcf67651bcf66520bef66520aef56552ccf56512ccf;
assign testcases[897] = 512'h10000fef10000fff97310adf92100dff80210eff70110aff70521ccf70522bbf10000fff00000fff76762bbf77661bbf76520aef766209ef67662cbf66613cbf;
assign testcases[898] = 512'h10000fef10000fff974109dfa2100dff80210eff80110aff80521bbf80522bbf10000fff00000fff76773abf78762abf77520aef766209ef67662cbf67623cbf;
assign testcases[899] = 512'h10000fef10000fffa84109dfa2100dff80210eff80110aef80531bbf80532bbf10000fff00000fff86873abf88762abf776209ef876209ef67772bbf67623bbf;
assign testcases[900] = 512'h10000fef10000fffa84108dfa2110cff90210dff902109ef80631abf80632abf10000fff00000fff878739af898729af876209ef877208ef78772bbf68723bbf;
assign testcases[901] = 512'h00000fff10000fff51100fff50000fff30000fff30000fff40100fef40100fef00000fff00000fff31110fef31110fef22100fff22100fff21110fef21100fef;
assign testcases[902] = 512'h00000fff10000fff52100fff61000fff30100fff40000fff40110fef40110fef00000fff00000fff32211fef32210fef32210fff32210eff32210fef32201fef;
assign testcases[903] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff50210fef50210fdf00000fff00000fff42221eef43220eef33210eff33210eff33221fdf33201fdf;
assign testcases[904] = 512'h00000fff10000fff63100eff61000fff40100fff40100eff50210edf50211edf00000fff00000fff43321eef43321eef43310eff43310dff33221edf33311edf;
assign testcases[905] = 512'h10000fff10000fff63200def71000fff50100fff50100dff50211edf50211edf00000fff00000fff43331edf44331edf43310dff43310dff34321edf33311edf;
assign testcases[906] = 512'h10000fef10000fff74210def71100eff50110fff50100dff60311ddf60311ddf00000fff00000fff54441ddf55431ddf54310dff54410cff44431edf44411edf;
assign testcases[907] = 512'h10000fef10000fff75210cef81100eff60110fff60110cff60421dcf60321dcf00000fff00000fff64542ccf55541cdf55410cff55510bff45441dcf45412dcf;
assign testcases[908] = 512'h10000fef10000fff86310bef82100eff70110eff60110bff70421ccf70421ccf00000fff00000fff65652ccf66551ccf65410bff65510bff56552dcf55512dcf;
assign testcases[909] = 512'h10000fef10000fff86310aef92100eff70210eff70110bff70421ccf70421ccf10000fff00000fff75762bcf67651bcf66520bef66520aef56552ccf56512ccf;
assign testcases[910] = 512'h10000fef10000fff97310adf92100dff80210eff70110aff70521ccf70522bbf10000fff00000fff76762bbf77762bbf76520aef766209ef67662cbf66623cbf;
assign testcases[911] = 512'h10000fef10000fff974109dfa2100dff80210eff80110aff80531bbf80522bbf10000fff00000fff76873abf78762abf77520aef766209ef67662cbf67623cbf;
assign testcases[912] = 512'h10000fef10000fffa84109dfa2100dff80210eff80210aef80631bbf80532bbf10000fff00000fff87873abf88762abf776209ef877208ef68772bbf67723bbf;
assign testcases[913] = 512'h10000fef10000fffa84108dfa2110dff90210eff802109ef80631abf80632abf10000fff00000fff878739af898729bf876209ef877208ef78772bbf68723bbf;
assign testcases[914] = 512'h30221edf30310def52100fff61000fff40100fff50100eff40100fef40100fef31321def31321ddf32110fef32110fef43310dff43310dff32110fef32100fef;
assign testcases[915] = 512'h30221edf30310def52100fff61000fff50100fff50100eff40100fef40100fef31321def31321ddf32110fef32110fef43310dff43310dff32110fef32100fdf;
assign testcases[916] = 512'h30221edf30310def52100fff61000fff50100fff50100eff40100fef50100fef31321def31321ddf32110fef32110fef43310dff43310dff32110fdf32200fdf;
assign testcases[917] = 512'h30221edf30310def52100fff61000fff50100fff50100eff40100fef50100fef31321def31321ddf32210fef32110fef43310dff43310dff32110fdf32200fdf;
assign testcases[918] = 512'h30331edf40320def51000fff50000fff40100fff40100eff40100fef40100fef41456cdf31335dde21110fef31111fef42310dff42310dff21110fef31101fef;
assign testcases[919] = 512'h30331edf40420def52000fff50000fff40100fff40100eff40100fef40100fef51442cdf41332ddf31110fef32110fef43310dff43310dff32110fef32100fef;
assign testcases[920] = 512'h30331edf40420def52000fff50000fff40100fff40100eff40100fef40100fef51442cdf41332ddf31110fef32110fef43310dff43310dff32110fef32100fef;
assign testcases[921] = 512'h30332edf40431def52000fff50000fff40100fff40100eff40100fef40101fef51445cdf41334ddf31110fef32111fef43310eff43310dff32111fef32101fef;
assign testcases[922] = 512'h30331edf40420def52000fff50000fff40100fff40100eff40100fef40100fef51542cdf41332dde31110fef32110fef43310dff43310dff32110fef32100fef;
assign testcases[923] = 512'h10000fef10000fff934109dfa1110dff80210eff80210aff80632bbf80632bbf00000fff00000fff73862bbf73762abf74620aef847209ef63662ccf63623cbf;
assign testcases[924] = 512'h10000fef10000fffa34109dfa1110dff80210eff80210aff80632bbf80632bbf00000fff00000fff73873abf73772abf74620aef847309ef63662ccf63723cbf;
assign testcases[925] = 512'h10000fef10000fff8c310cef83100eff90210eff902109ef60421dcf60421dcf00000fff00000fff5c552cdf5c551ddf858319ef96a418ef4b441dcf4b512dcf;
assign testcases[926] = 512'h10000fef10000fff73310cef81100eff90210eff902109ef60421dcf60421dcf00000fff00000fff53542cdf53551ddf848319ef949417ef43441dcf43412dcf;
assign testcases[927] = 512'h10000fef10000fff85310bef81100eff90320eff90210aef70531ccf70422ccf00000fff00000fff64652ccf55552ccf858319ef96a418ef45552dcf55513dcf;
assign testcases[928] = 512'h10000fef10000fff83310bef81100eff90210eff902109ef70421ccf70421ccf00000fff00000fff63552ccf54551ccf858319ef959317ef43452dcf53512dcf;
assign testcases[929] = 512'h10000fef10000fff8f310cef84100eff90210eff90210aef60421dcf60421dcf00000fff00000fff5f552ddf5f551ddf868319ef96a418ef4f441ddf4f512dcf;
assign testcases[930] = 512'h10000fef10000fff73310cef81100eff90210eff802109ef60421dcf60421dcf00000fff00000fff53542cdf53541ddf848319ef949317ef43441dcf43412dcf;
assign testcases[931] = 512'h10000fef10000fff86310bef92100eff90210eff80210aef70532ccf70422ccf00000fff00000fff65662ccf66662ccf858319ef959418ef56562dcf56623dcf;
assign testcases[932] = 512'h10000fef10100fffb76206bdc2210cffc0420cffc03215efa095299da084399d10000fff00000fff96ba489d97a9389ec7c414dfd7f512df76993aad76a35a9d;
assign testcases[933] = 512'h10000fef10000fffb45106cfb1110cffc0320dffb03106ef907429afa07429af00000fff00000fff93a938af849828afc5a415efc5c413df73783bbf74824aaf;
assign testcases[934] = 512'h10000fef10000fffb65107dfb2110cffc0321dffc03116efa07429afa07329af01001fff01001fff959839af968829afcbb415efdad414df76772bbf76824aaf;
assign testcases[935] = 512'h10000fef10000fff84310bef81100eff80210eff80210aff70531ccf70422ccf00000fff00000fff63652ccf64651ccf84731aef848318ef53552dcf53513dcf;
assign testcases[936] = 512'h10000fff10000fff84310bef91100eff80210eff80210aff70531ccf70522ccf00000fff00000fff64652ccf64651ccf85731aef858318ef54552dcf54513dcf;
assign testcases[937] = 512'h10000fef10000fff85310bef91100eff80210eff80210aff70532ccf70532ccf00000fff00000fff65762ccf66662ccf85831aef859418ef55562dcf55623dcf;
assign testcases[938] = 512'h00000fff10000fff87310cef82100eff70210eff70210bff60421dcf60421dcf00000fff00000fff57552cdf56551ddf74621aef747319ef46442dcf46512dcf;
assign testcases[939] = 512'h10000fef10000fff85410bef91110eff80210eff80210aff70532ccf70532ccf00000fff00000fff64773ccf65662ccf85731aef859319ef55562dcf55623dcf;
assign testcases[940] = 512'h10000fef10000fff85310bef91100eff80210eff80210bff70532ccf70532ccf00000fff00000fff65763ccf66662ccf75731aef858319ef55562dcf55623dcf;
assign testcases[941] = 512'h10000fff10000fff95410aef91110eff80210eff80210aff70532ccf70532ccf00000fff00000fff64773bcf65662ccf85731aef859319ef55562dcf55623dcf;
assign testcases[942] = 512'h10000fff10000fff95410aef91100eff80210eff80210aff70531ccf70532ccf00000fff00000fff64763bcf65662ccf74731aef848319ef54562dcf54623dcf;
assign testcases[943] = 512'h41331cce50420cdf86410bef82110effc0310dffc02107ef80742bbf80732bbf55442bdf55442cce66983ccf67872bcfcaa315efcab314ef68783cbf68824bbf;
assign testcases[944] = 512'h40451cce50531bdf86210bef81100effb0310dffc02107ef80421bbf80421bbf55552bdf55553bce65441bcf66541bcfc9a315efc9a314ef66541bbf76612bbf;
assign testcases[945] = 512'h30551dde30531def74210cef71100eff90310eff902109ef70421ccf70421ccf33563cdf33563dde54431ddf54541ccfa79317efa7a316ef55541ccf55612cbf;
assign testcases[946] = 512'h31441ddf40430cef74210cef81100effa0310effa02109ef70421ccf70421ccf34442ddf34442dde54442ddf55441cdfa6a418efa6a417ef55452dcf55513ccf;
assign testcases[947] = 512'h31441dde40430cef84210cef81100effa0320effa02108ef80521ccf80422ccf34442cdf35442dde64552ccf65551ccfb6a417efb6b416ef55552ccf65623ccf;
assign testcases[948] = 512'h31341dde41420def78210def72100fffa0221effa02119ef70421dcf70322dcf36442ddf37342dde67442ddf6a442cdfa89428efa8a417ef5a542dcf6b513ccf;
assign testcases[949] = 512'h31331edf30320def74210cef81100eff90221eff90211aff70421ccf70422ccf35331def35332ede53442ddf54441ddf969419ef969419ef54552dcf55513dcf;
assign testcases[950] = 512'h31332edf30320def73210cef81100eff90221eff90211aff70421ccf70421ccf34333def34333ede53442ddf53451ddf959419ef959318ef54542dcf53513dcf;
assign testcases[951] = 512'h20220eef20210eef62200eff71000fff70211fff70211cff60321ddf60321ddf23221eef23221eef42332edf42331edf74731bff74731aff43342edf42413edf;
assign testcases[952] = 512'h20220eef20210eff62100eff61000fff60210fff70110cff50311edf50211edf23221eef23221eef42331eef43331eef74731bff74731bff43331edf43412edf;
assign testcases[953] = 512'h40551cce50531bde84210bef91100effb0310dffb02107ef80521bbf80521bbf44552cde44553cce75652bcf76651bcfc7b415efc7b414ef76652bbf76723baf;
assign testcases[954] = 512'h10000fff10000fff94410aef91100eff80210eff80210aff70531ccf70532ccf00000fff00000fff74763bcf64662ccf74731aef848319ef54562dcf54623ccf;
assign testcases[955] = 512'h10000fff10000fff95410aef91110eff80210eff80210aff70632ccf70532ccf00000fff00000fff65773bcf66672ccf75731aef858319ef55672dcf55624ccf;
assign testcases[956] = 512'h00000fff10000fff74310cef81100eff60210fff60110cff60421ddf60422ddf00000fff00000fff53652ddf54551ddf63631cff64731bff43452edf43513edf;
assign testcases[957] = 512'h10000fef10000fffa75109dfa2110dff90210eff902109ef90742abf90643abf00000fff00000fff86994abf87882abf968318efa6a317ef66783cbf76824bbf;
assign testcases[958] = 512'h41451cce40531cdf95310adf91100dffc0321dffc03217ef90632abf90632abf47452cdf47443cce84763abf76762abfc8c516efc8c515ef76772bbf86824baf;
assign testcases[959] = 512'h10110fef10100fff71310def80100eff90210effa02109ef60411edf60411edf10000fff10000fff41431edf51531ddfa58208efb5a205ef31321edf41311edf;
assign testcases[960] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58208efc5a205ef31321edf41311edf;
assign testcases[961] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58208efc5a205ef31321edf41311edf;
assign testcases[962] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58208efc5a205ef31321edf41311edf;
assign testcases[963] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc6a205ef31321edf41311edf;
assign testcases[964] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[965] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[966] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[967] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[968] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[969] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[970] = 512'h10110fef10100fff82310def90100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[971] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[972] = 512'h10110fef10100fff82310def90100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[973] = 512'h10110fef10100fff82310def90100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc6a205ef31321edf41311edf;
assign testcases[974] = 512'h10110fef10100fff82310def90100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc6a205ef31321edf41311edf;
assign testcases[975] = 512'h10110fef10100fff82310def90100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[976] = 512'h10110fef10100fff82310def90100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc6a205ef31321edf41311edf;
assign testcases[977] = 512'h10110fef10100fff82310def90100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc6a205ef31321edf41311edf;
assign testcases[978] = 512'h10110fef10100fff82310def80100eff90210effa02109ef60411edf60411ddf10000fff10000fff41431edf51531ddfa58207efc5a205ef31321edf41311edf;
assign testcases[979] = 512'h10000fef10100fff82310def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321eef51431edf947209efa49207ef31321fdf31311edf;
assign testcases[980] = 512'h10000fef10100fff82310def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431edf948209efa49207ef31321edf31311edf;
assign testcases[981] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431edf948209efb49207ef31321edf31311edf;
assign testcases[982] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431ddf948209efa49207ef31321edf31311edf;
assign testcases[983] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431ddf948209efb49207ef31321fdf31311edf;
assign testcases[984] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431ddf948209efb49207ef31321edf31311edf;
assign testcases[985] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431edf948209efb59207ef31321edf31311edf;
assign testcases[986] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431ddf948209efb49207ef31321edf31311edf;
assign testcases[987] = 512'h10000fef10100fff82310def80100fff80210eff90210aef60411edf60311edf10000fff10000fff41321edf51431ddf948209efb59207ef31321edf31311edf;
assign testcases[988] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431ddf948209efb59206ef31321edf31311edf;
assign testcases[989] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321eef51431ddf948209efb59207ef31321edf31311edf;
assign testcases[990] = 512'h10000fef10100fff82210def80100fff80210eff90210aef60311edf60311edf10000fff10000fff41321edf51431ddf948209efb59206ef31321edf31311edf;
assign testcases[991] = 512'h10000fef10100fff82210def80100fff80210eff90210aef60311edf60311edf10000fff10000fff41321edf51431ddf948209efb59206ef31321edf31311edf;
assign testcases[992] = 512'h10000fef10100fff82210def80100fff80210eff90210aef60311edf60311edf10000fff10000fff41321edf51431ddf948208efb59206ef31321edf31311edf;
assign testcases[993] = 512'h10000fef10100fff71210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431ddf948209efb49207ef31321edf31311edf;
assign testcases[994] = 512'h10000fef10100fff72210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431ddf948209efb59207ef31321edf31311edf;
assign testcases[995] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321eef51431ddf948209efb59206ef31321edf31311edf;
assign testcases[996] = 512'h10000fef10100fff82210def80100fff80210eff90210aff60311edf60311edf10000fff10000fff41321edf51431ddf948208efb59206ef31321edf31311edf;
assign testcases[997] = 512'h10000fef10100fff72210def80100fff80210eff90210aef60311edf60311edf10000fff10000fff41321edf51431ddf948209efb59207ef31321edf31311edf;
assign testcases[998] = 512'h10000fef10100fff72210def80100fff80210eff90210aef60311edf60311edf10000fff10000fff41321edf51431ddf948209efb59206ef31321edf31311edf;
assign testcases[999] = 512'h10000fef10100fff71200eff80100fff70210fff80100bff60310edf60311edf00000fff00000fff41321eef51321eef83610aef947109ef31210fdf31201fdf;


  
  localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
  wire [$clog2(CLASS_CNT)-1:0] prediction;

  // Instantiate module under test
 gasId_bnn1_bnnseq #() dut (
    .features(sample),
    .clk(clk),
    .rst(rst),
    .prediction(prediction)
  );
  
  always #halfPeriod clk <= ~clk;

  integer i;
  initial begin
    $write("["); //"
    for(i=0;i<TEST_CNT;i=i+1)
        runtestcase(i);
    $display("]");
    $finish;
  end

  localparam [$clog2(CLASS_CNT)-1:0] maxclass = CLASS_CNT-1;

  task runtestcase(input integer i); begin
    sample <= testcases[i];
    rst <= 1;
    clk <= 0;
    #period
    rst <= 0;
    #period
    #((FEAT_CNT+HIDDEN_CNT-1)*period)
    $write("%d, ",(maxclass-prediction));
  end
  endtask

endmodule
