
















module gasId_tnn1_tnnpaarter #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 37488'h00540364000102ce03630001035a03620001034f036100010333036000010352035f00010346035e000102b9035c00010345035b0001030603590001035703580001031e03560001031003550001030f0354000102da035100010319035000010314034d00010324034c0001030a0349000102520348000103380347000102c20343000102b00342000103160341000102cb034000010330033f0001032d033e0001032f033c0001031c033b000102bc0339000103250337000102f10334000102fa033100010309032e0001032a032c000102bd032900010320032800010323032600010308031d00010304030c0001034b035d00000344035300000321034e00000327034a00000305033d000002fb033a0000031303360000030b0335000003000332000002fc032b000002db0322000002d4031f000002f8031b000002e8031a000002d10318000002d90317000002f00315000003030312000002a90311000002c8030e000002d3030d000002fd0307000002e303020000029c0301000002ca02ff000002ec02fe000002d702f9000002c002f70000027802f60000029d02f5000002b802f40000028b02f3000002c702f20000028102ef0000028302ee0000029402ed0000027c02eb0000026d02ea0000025402e9000002be02e70000029902e6000002b402e5000002b602e40000028602e2000002ac02e10000027502e0000002cc02df000002cd02de0000029f02dd0000028402dc0000029202d80000024802d6000002a102d50000025802d20000024a02d0000002a802cf0000024002c90000028a02c60000026f02c50000028e02c40000025d02c30000029a02c10000028502bf0000022002bb0000026102ba0000024e02b70000027902b50000027f02b30000021502b20000024f02b10000020a02af0000020f02ae0000021602ad0000027702ab0000027202aa000001f602a70000024b02a60000024c02a50000025c02a40000026602a30000025102a20000027e02a000000280029e00000287029b000001d002980000026502970000027d02960000022802950000021c02930000027b0291000002730290000001ee028f00000212028d00000270028c000001d402890000025602880000019602820000026e027a000002430276000001e402740000026b027100000247026c0000025e026a000001fd02690000024402680000024102670000019502640000023902630000023f026200000233026000000188025f00000224025b0000020c025a000001e20259000002380257000001b30255000001cd025300000205025000000229024d000001e80249000002370246000001b10245000001c30242000001da023e00000235023d00000226023c00000223023b00000202023a000002110236000002040234000001a402320000020702310000017902300000022c022f0000021b022e000001dd022d000001e3022b00000200022a000001b80227000001cb02250000020e02220000020102210000018a021f000001db021e000001de021d000001ac021a000001f40219000001ef0218000001720217000001ec0214000001d30213000001dc0210000001f0020d0000016a020b000001fb0209000001bc0208000001f20206000001c50203000001c201ff000001e501fe000001c601fc0000016d01fa0000014e01f9000001bd01f8000001e901f7000001af01f5000001bb01f30000014901f1000000c201ed0000010f01eb000001c101ea0000011f01e70000015c01e60000019d01e1000001a601e0000001ca01df0000015d01d9000001a001d8000001a901d70000017401d6000000ad01d50000013f01d20000012f01d10000018701cf0000013c01ce0000017001cc000001a201c9000001bf01c80000016401c70000019101c40000016901c00000014101be0000015d01ba0000016501b90000019e01b70000012f01b60000018901b50000016001b40000018501b20000016e01b00000017601ae0000018c01ad0000018401ab0000014f01aa0000014401a80000017c01a70000018601a50000011501a30000016901a100000121019f00000174019c00000192019b0000017a019a0000013d01990000015e0198000000f401970000018e01940000017501930000017f019000000144018f00000173018d00000181018b0000013301830000011101820000015101800000015a017e00000160017d00000168017b0000017701790000017601780000016a01780000017301750000013501720000016b017100000162017100000162017000000163016f00000158016f00000132016e00000143016c000000f9016c000000c00168000001520167000001650166000001630166000000fe01640000015f016100000137016100000130015f00000156015e00000159015a000000f501580000013401560000014701550000014101550000009101540000005a0154000001280151000001280150000000ba01500000012e014f000000a2014e00000143014b00000138014a000000f5014a0000010d01490000013e01470000012201460000011e0146000001240140000001230140000000ab013f0000011f013e00000080013d000000e5013c00000079013a0000013001390000012401390000011a0138000000fb0137000000f90136000000fc0135000000e40134000000e60133000000f601310000012a012e00000116012b000000e80127000000d101270000010e0126000000810126000001140123000000d20121000000c8011e00000115011c0000010f011c00000108011a000001120117000000e50117000000fd01160000010c01120000010b011100000105010e000000be010d00000106010b000000ca010a00000088010a000000ed0106000000fa0105000001010104000000f10104000000cb00fe000000df00fc000000cf00fa000000c100fa000000c500f9000000ee00f8000000a200f7000000e300f4000000d700f4000000cc00f30000008e00f2000000e900f0000000d900ef000000b200ed0000005600ed000000b400ec000000ac00eb000000cc00e7000000e400e6000000bd00e6000000cd00e5000000c100e40000008300e3000000b800e2000000ad00e1000000c100e00000009500e00000008200e0000000c600dd000000ab00dc0000008a00db000000d800da000000b100d6000000be00d50000009200d3000000a200d2000000c400d1000000b400cf000000c900ce000000b900c9000000a400c8000000af00c7000000c500c6000000b600c4000000b800bf000000aa00bf000000ad00bd000000a100bd0000003700bd000000b600bc0000002900bc0000009a00bb0000007d00b8000000af00b7000000b200b6000000b000b50000005c00b50000004200b50000009800b1000000a600b00000002600af0000007c00ae0000008100ad0000007800ac0000007200a90000009100a80000000200a80000009400a50000008200a20000003c00a10000000c00a10000006200a00000009b009f00000068009f0000003e009f00000048009e0000008c009d0000007d009b0000008300990000009000970000008800960000007900920000007800920000004200920000003d00910000003f00900000006e008e00000010008a0000004500890000002200890000004800870000006500860000004c00860000005200850000002c00850000005f008200000068007e00000067007e00000073007c00000033007b00000055007a0000007200780000006c00770000006000760000005a00760000006500740000002300740000001600730000006d00710000001c00710000006c00700000004b00700000005d006f00000009006e00000042006d00000017006d0000001400640000002100620000005a006100000021006000000059005f00000001005b00000000005a0000005300580000003d00550000000a00520000002a00510000000e00500000000b004f00000049004e0000002e004c00000003004a0000000d00490000000500460000001b00450000003600440000003400410000001c004100000031004000000020003c00000028003b0000002500380000000400380000002200360000002000360000000d00320000002600300000001b002d00000003002c00000004002b00000019002a0000001900230000000c001f00000010001e00000018001a0000000500160000000800120000000200070000000300040000010c01770001012b016b0001015201670001014b0159000100700136000100560131000100e30108000100aa00c100010020009d0001006e016d00000101015c00000068013a00000033013200000071012a0000000201220000006c0114000000f500fd0000004a00cd0000001000af0000004200a80000006e009a0000006200f700010066015b0001001f015700010109015300010096014d000100f6014800010004012d000100e7012c000100d001200001007f011d0001004b01130001000f01000001008d00e90001009400e20001002400e10001008f00dd000100d000d80001006100d60001006b00d30001000600b1000100a500a800010095009800010063008d0001001d008000010014003a00010107014c000000f80145000000c90142000000f0013b000000da01290000008c01250000008a011b000000f20119000000c40118000000dc0110000000b30103000000d901020000003200ff0000003100fb000000db00f30000005500f1000000cf00ef0000003500ee0000009e00ec000000c800eb0000009700e80000002d00df0000008400d70000007000d20000005000cd000000c300cc0000000000c50000003900c30000009800bf0000006900be0000008100bb0000000800bb0000006b00b7000000a700b40000001300b40000008400b20000009f00b00000007300ac0000004000aa0000007a00a90000009e00a7000000a300a40000002100a00000005c009b0000002a009b0000002c009900000046008f00000087008e00000081008c00000038008800000028008600000082008500000069008500000035007e00000041007c0000002c00770000004700760000003400740000004b006f0000001e006e00000008006d00000060006a0000006500680000001a00600000003d005d0000003800580000000400580000001300570000005200540000002b005100000009005000000014004e0000000d004d0000004100490000002900490000004500480000000300470000002d004000000017003f00000012003c00000034003b00000022003900000028003200000011002e0000000200270000000e00150000007400d10001005300b70001001200ab00010041008e0001003000510001002900510001001b004500010011003c0001005f00d50000007800c60000004d00b80000002c00a90000007300990000003f0095000000390057000000ce00ea0001005200de0001002a00cb0001001000ca000100b100b50001005400a200010015007c0001000b007b0001003d00590001003100560001007d00d40000008000c20000003000c00000008900bc0000009d00b60000000c00b20000007800a70000001a00a50000006500a000000062009f00000070009e0000008300980000007200970000006a009100000019009000000018008f00000020008b0000000e00850000002f007f0000005b006100000042004300000036003e0000001c003500000017002d0000001d002200000019001b00000012008a0001006900790001000500160001000f00c7000000020048000000b900ba00010013009c0001004f005e00010033005a0001000400b30000008c00b00000000c00af0000002300a60000002000930000003b007b00000032006d0000003a006700000025005c0000000100440000002100310000000700240000008200a700010009008b0001000100530001002b004e00010010006800000014001c000000a900ad0001000200ac0000007800ab000000a800aa0000002400a2000000450074000000a500a60001002c009f00000030009e0000002000980001004100a000000072007a0000009b00ae00000018005a0000002800a400010054009900010001009d00000034005800010010003c000100a100a300010097009c00000069009500010014008c00000003001200010091009a00000059008f0000006000680000008b00960000000400090000001b008a0000003b00940001009200930000008e00900000005b007900000071007300000050008500010041005c00000074007c00000052008d0001006100700001008200890001004200880000000000860000003300530000004a00870000001100190000004b008300000051006a0001001c00840000002a00620000001300810000007b00800001001a00430001002300490000004000440000000c002200010048004c00000063006b00000008002b00010064006c0000000a000b0000 ;
localparam YMAP = 1280'h0000036d000103660000036c000103750001037000000378000103870000037e000103650000038c0000038b000103740000036a00000383000103770000036b0001038500000384000103730000037c0001036900000386000003710001036700010382000003810000037d00010368000003800001037b0000036e0000037a0000038800010389000003720000036f000103760001038a000003790001037f;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 240'b000100000000000000010000000000000000000010000000000000010100000000010001000100000000000000100000000000000000000000000000000000010011010000000000000000000000000000100000000100000010000100100001000000000000010000100000000010000000010100000000 ;
localparam WNNZ = 240'b000100000000001001110010001000000101100010010000000000010110000000010001001100000000000000100000000000100001000000000000000011010011011000000010000100100100000100100000100100000010100100101111000000011000010110100100010010000100010100000100;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
wire [SUM_BITS-1:0] scorarr [CLASS_CNT-1:0];
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;

generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam adsub = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(adsub)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] <= 0;
end
endgenerate

function [7:0] zerocnt(input integer k);
    integer i,j;
    reg [HIDDEN_CNT-1:0] neur1;
    begin
        i = 0;
        neur1 = WNNZ[k*HIDDEN_CNT+:HIDDEN_CNT];
        for(j=0;j<HIDDEN_CNT;j=j+1)
            i = i + !(neur1[j]);
        zerocnt = i;
    end
endfunction

function [7:0] minzc(input integer k);
    integer i,j,h;
    begin
        i = HIDDEN_CNT;
        for(j=0;j<CLASS_CNT;j=j+1) begin
            h = zerocnt(j);
            if(h<i)
                i = h;
        end
        minzc = i;
    end
endfunction

localparam MINZC = minzc(0);

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    localparam Wuse = WNNZ[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wuse[j]) begin
            if(Wneur[j])
                tmpscore = tmpscore + hidden[j];
            else 
                tmpscore = tmpscore + hidden_n[j];
        end
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = 2*tmpscore + zerocnt(i) - MINZC;
    /* assign scorarr[i] = 2*tmpscore + zerocnt(i) - MINZC; */
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
