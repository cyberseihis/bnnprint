`timescale 1us/1ns









module tbcardio_bnn1_bnnseq #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000


)();

  
  reg [FEAT_BITS*FEAT_CNT-1:0] sample;
  wire [FEAT_BITS*FEAT_CNT-1:0] testcases [TEST_CNT-1:0];
  reg rst;
  reg clk;
  parameter Nsperiod=50000;
  localparam period=Nsperiod/500;
  localparam halfPeriod=period/2;


assign testcases[0] = 76'h46980212600181d0004;
assign testcases[1] = 76'h199a25a3b0230413028;
assign testcases[2] = 76'h199a24a3b0240413018;
assign testcases[3] = 76'h199a0a70a0270514018;
assign testcases[4] = 76'h199a0870a0060513028;
assign testcases[5] = 76'ha45254b0d8900d37018;
assign testcases[6] = 76'hd45155b0d8600e46018;
assign testcases[7] = 76'h07780012600511f0005;
assign testcases[8] = 76'h07780012600411f1005;
assign testcases[9] = 76'h07780112600310f2005;
assign testcases[10] = 76'h1bbb0291b01924b100d;
assign testcases[11] = 76'h1bbb0491b01914b100d;
assign testcases[12] = 76'h0999044660240334227;
assign testcases[13] = 76'h199a025380120333447;
assign testcases[14] = 76'h598a067294620523e47;
assign testcases[15] = 76'h3889037294330512827;
assign testcases[16] = 76'h498a0480b0330432827;
assign testcases[17] = 76'h3889047294340511717;
assign testcases[18] = 76'h2879055194330423917;
assign testcases[19] = 76'h28892582a4520444f47;
assign testcases[20] = 76'h86590c81bc230443907;
assign testcases[21] = 76'h288908a1c4220431827;
assign testcases[22] = 76'h94422ab1d8210551607;
assign testcases[23] = 76'h07780019100201f0007;
assign testcases[24] = 76'h088900191001e0f1007;
assign testcases[25] = 76'h0778011a1001d0f0005;
assign testcases[26] = 76'h0788013b200220f0005;
assign testcases[27] = 76'h0778001a1001c0f0005;
assign testcases[28] = 76'h487926a0c4a30a41508;
assign testcases[29] = 76'h566909a0d0820e30208;
assign testcases[30] = 76'h377908b0d0c40a31408;
assign testcases[31] = 76'h466809b0d0a20f22208;
assign testcases[32] = 76'h28792aa0d0750641208;
assign testcases[33] = 76'h17780c81b0170831364;
assign testcases[34] = 76'h17892880b0140731244;
assign testcases[35] = 76'h17780aa0d0080834334;
assign testcases[36] = 76'h16670880b0360824343;
assign testcases[37] = 76'h16670790c0250732022;
assign testcases[38] = 76'h16670790c0160822133;
assign testcases[39] = 76'h16770680b0040533263;
assign testcases[40] = 76'h1677264190140536262;
assign testcases[41] = 76'h16770581b0040534122;
assign testcases[42] = 76'h1778054180040362113;
assign testcases[43] = 76'h17782ca0d0040463023;
assign testcases[44] = 76'h166706b0d0450a21005;
assign testcases[45] = 76'h166707b0d0450b21005;
assign testcases[46] = 76'h17780ca0d0270b13005;
assign testcases[47] = 76'h27780aa0d0270b23015;
assign testcases[48] = 76'h477906b0d0450f23015;
assign testcases[49] = 76'h1eee06a4b015043604f;
assign testcases[50] = 76'h1eee04ae5004034402f;
assign testcases[51] = 76'h4bab26b0d057097600f;
assign testcases[52] = 76'h699707b0d4610c5600f;
assign testcases[53] = 76'h0bcc025c301271a000d;
assign testcases[54] = 76'h0bbb034d1002c0c000c;
assign testcases[55] = 76'h0bbb2b91b02492a000d;
assign testcases[56] = 76'h0bbb2b91b01493a000d;
assign testcases[57] = 76'h0ccc016e1002716300c;
assign testcases[58] = 76'h0bcc016e2002516300c;
assign testcases[59] = 76'h0bcb04849002024303b;
assign testcases[60] = 76'h0bcc048c4002326302c;
assign testcases[61] = 76'h0bcc027e2002416202c;
assign testcases[62] = 76'h0abb005c2004033100b;
assign testcases[63] = 76'h09aa0a94a0040333019;
assign testcases[64] = 76'h0aaa09849004033301a;
assign testcases[65] = 76'h0bcc015e1002716200d;
assign testcases[66] = 76'h0ccd388590044272019;
assign testcases[67] = 76'h0bcc028a5003025203a;
assign testcases[68] = 76'h0bcc028a5003025203a;
assign testcases[69] = 76'h0ccd046c3004017400b;
assign testcases[70] = 76'h0ccd036d2004017301b;
assign testcases[71] = 76'h1abb00739005039206a;
assign testcases[72] = 76'h1abb02739004039004a;
assign testcases[73] = 76'h1abb02739006049305a;
assign testcases[74] = 76'h1bbc03739005039507a;
assign testcases[75] = 76'h0ccc0264800402b100e;
assign testcases[76] = 76'h0bcc006d200312a100d;
assign testcases[77] = 76'h1bbb2371a004035102c;
assign testcases[78] = 76'h1bbb2571a007045101c;
assign testcases[79] = 76'h1bbb04a1c007045202c;
assign testcases[80] = 76'h1bbb2461a008045100c;
assign testcases[81] = 76'h0bbb28a1c006036101c;
assign testcases[82] = 76'h0bbb27a1c005026100c;
assign testcases[83] = 76'h1ccc0472a000037104c;
assign testcases[84] = 76'h1ddd0492b004026116c;
assign testcases[85] = 76'h1ddd0493a000026117c;
assign testcases[86] = 76'h1bbc0460a007046103c;
assign testcases[87] = 76'h09990490c014036010a;
assign testcases[88] = 76'h0abb0493a00451b000a;
assign testcases[89] = 76'h3a9b6bb0d022058001a;
assign testcases[90] = 76'h1ccd016c200250b101a;
assign testcases[91] = 76'h0bbb044d1002c0c000c;
assign testcases[92] = 76'h0bbb024d1002c0c000c;
assign testcases[93] = 76'h0bbb034b2001d0c000c;
assign testcases[94] = 76'h0bbb004d1001d0d100c;
assign testcases[95] = 76'h0bbb015c200311a000c;
assign testcases[96] = 76'h0bbb235a300350b000c;
assign testcases[97] = 76'h0bcc0354701291a000c;
assign testcases[98] = 76'h0bcc025c301271a000c;
assign testcases[99] = 76'h089927a780020411046;
assign testcases[100] = 76'h1889036380241431026;
assign testcases[101] = 76'h0889354750150331046;
assign testcases[102] = 76'h0899044370050331036;
assign testcases[103] = 76'h0889003a20030240016;
assign testcases[104] = 76'h0889244370050420016;
assign testcases[105] = 76'h17782491b0550622136;
assign testcases[106] = 76'h166826a0d0440920106;
assign testcases[107] = 76'h1788078390140422026;
assign testcases[108] = 76'h178827a2c0420523136;
assign testcases[109] = 76'h0788243450060330006;
assign testcases[110] = 76'h178909b4b0410521126;
assign testcases[111] = 76'h099a09a4a0040451047;
assign testcases[112] = 76'h099a05a780030352027;
assign testcases[113] = 76'h0899246950040261007;
assign testcases[114] = 76'h587a2ca0d0800c24037;
assign testcases[115] = 76'h46693690c0700b22007;
assign testcases[116] = 76'h755827a0d4160a32005;
assign testcases[117] = 76'h0778034750520243025;
assign testcases[118] = 76'h0778034650410242015;
assign testcases[119] = 76'h0778034650310332015;
assign testcases[120] = 76'h17793c91b0525274005;
assign testcases[121] = 76'h0778066480316182005;
assign testcases[122] = 76'h1778273170413272005;
assign testcases[123] = 76'h277928b2c0210342025;
assign testcases[124] = 76'h1667232274310333005;
assign testcases[125] = 76'h0ddd0075800330b300f;
assign testcases[126] = 76'h0ddd006f100240c200f;
assign testcases[127] = 76'h0ddd0075800411b100f;
assign testcases[128] = 76'h0ddd006f100220b100f;
assign testcases[129] = 76'h0ddd03748003619000f;
assign testcases[130] = 76'h0ddd007f1002719000f;
assign testcases[131] = 76'h0ddd01648003519000f;
assign testcases[132] = 76'h0ded007f1001a1a000f;
assign testcases[133] = 76'h0ddd048c400310a701f;
assign testcases[134] = 76'h0ddd048c400201a401f;
assign testcases[135] = 76'h0ddd007f200320c400f;
assign testcases[136] = 76'h0ddd048c400201a401f;
assign testcases[137] = 76'h0ddd007e200230c300f;
assign testcases[138] = 76'h0eed009e300311a601f;
assign testcases[139] = 76'h0efd029e400321a401f;
assign testcases[140] = 76'h0dee018f200301a100f;
assign testcases[141] = 76'h2cccf9a0d018047102e;
assign testcases[142] = 76'h0ddd04868004028100e;
assign testcases[143] = 76'h1ccc87a0d00b047101e;
assign testcases[144] = 76'h1abb0981b005128204b;
assign testcases[145] = 76'h0bbb04839001028103b;
assign testcases[146] = 76'h0abb27739006228101b;
assign testcases[147] = 76'h0bcb04739006128201d;
assign testcases[148] = 76'h0bcc24748003228001d;
assign testcases[149] = 76'h0bcc266a4003319301c;
assign testcases[150] = 76'h0bcc046a400341a100c;
assign testcases[151] = 76'h0bcb045a4003219100c;
assign testcases[152] = 76'h2bbc2b70b013046304a;
assign testcases[153] = 76'h189803b970040343026;
assign testcases[154] = 76'h078804b970050252006;
assign testcases[155] = 76'h0788024930032263015;
assign testcases[156] = 76'h0788023920032163015;
assign testcases[157] = 76'h0788013a20032263015;
assign testcases[158] = 76'h0788013a30012255055;
assign testcases[159] = 76'h0788024a30011243035;
assign testcases[160] = 76'h0788014a30013253025;
assign testcases[161] = 76'h0788014a30012253025;
assign testcases[162] = 76'h0778024270132244025;
assign testcases[163] = 76'h0788224560032243025;
assign testcases[164] = 76'h0788043550032242025;
assign testcases[165] = 76'h199a0191b01d0791028;
assign testcases[166] = 76'h199a0191b00f0891018;
assign testcases[167] = 76'h099a02a1c00813c1018;
assign testcases[168] = 76'h099a05a3b00502c1018;
assign testcases[169] = 76'h0778042640027171013;
assign testcases[170] = 76'h0678051160124172003;
assign testcases[171] = 76'h0778011910025181003;
assign testcases[172] = 76'h0778236480130342014;
assign testcases[173] = 76'h0778336480040341014;
assign testcases[174] = 76'h0778056480041341014;
assign testcases[175] = 76'h078806a1c0030342024;
assign testcases[176] = 76'h0788044180040251004;
assign testcases[177] = 76'h199908a3b0130443054;
assign testcases[178] = 76'h0778033650140332014;
assign testcases[179] = 76'h199a0aa1c0020441044;
assign testcases[180] = 76'h188829a3b0050432024;
assign testcases[181] = 76'h4ccb3ab0d0010c53089;
assign testcases[182] = 76'h1778244180210450007;
assign testcases[183] = 76'h18892680b0530663008;
assign testcases[184] = 76'h8dc928b0d0120b41038;
assign testcases[185] = 76'h489935a0d0750856038;
assign testcases[186] = 76'h0999044280070481008;
assign testcases[187] = 76'h0ccd377c40044272019;
assign testcases[188] = 76'h1ccd377c40043273019;
assign testcases[189] = 76'h0bcc028a50030341029;
assign testcases[190] = 76'h0ccd378590044272009;
assign testcases[191] = 76'h0ccd046c3004017301b;
assign testcases[192] = 76'h0ccd039d4003118101b;
assign testcases[193] = 76'h0ccd036d3004017301b;
assign testcases[194] = 76'h0ccc026e1002319400d;
assign testcases[195] = 76'h0ccc026e1002219200d;
assign testcases[196] = 76'h0ccd036e200231a200d;
assign testcases[197] = 76'h0ccc006d2004118100c;
assign testcases[198] = 76'h0ccc017e2002018101c;
assign testcases[199] = 76'h0778052170141190004;
assign testcases[200] = 76'h0778042170050180004;
assign testcases[201] = 76'h0778022820032190004;
assign testcases[202] = 76'h0778202920032190004;
assign testcases[203] = 76'h07780029200301a0004;
assign testcases[204] = 76'h0778211920023180004;
assign testcases[205] = 76'h0778002a10022190004;
assign testcases[206] = 76'h0778042170050290004;
assign testcases[207] = 76'h0778031260050190004;
assign testcases[208] = 76'h0889043640020171025;
assign testcases[209] = 76'h08890029200201a0005;
assign testcases[210] = 76'h0899083550020181166;
assign testcases[211] = 76'h0899013b10020180016;
assign testcases[212] = 76'h08990771a0010281046;
assign testcases[213] = 76'h0899033370020170026;
assign testcases[214] = 76'h08990432700311a1016;
assign testcases[215] = 76'h09990349300301a1016;
assign testcases[216] = 76'h08890442800411b0006;
assign testcases[217] = 76'h08890442800411a0006;
assign testcases[218] = 76'h199a283270151291046;
assign testcases[219] = 76'h099a036290060190026;
assign testcases[220] = 76'h0899094370040190127;
assign testcases[221] = 76'h0899033a20020190007;
assign testcases[222] = 76'h0899055090050270017;
assign testcases[223] = 76'h0899025a30020270017;
assign testcases[224] = 76'h0999035b30020190017;
assign testcases[225] = 76'h0899033a20020190007;
assign testcases[226] = 76'h0899024270040280056;
assign testcases[227] = 76'h1898024270050280026;
assign testcases[228] = 76'h0899023270040270026;
assign testcases[229] = 76'h0889062080050190025;
assign testcases[230] = 76'h0889044560030190015;
assign testcases[231] = 76'h0889022260041180005;
assign testcases[232] = 76'h0889044560030190015;
assign testcases[233] = 76'h0889022260041180005;
assign testcases[234] = 76'h0889022260041180005;
assign testcases[235] = 76'h0888032270030190024;
assign testcases[236] = 76'h0788002a20030190014;
assign testcases[237] = 76'h0888002a200211a0024;
assign testcases[238] = 76'h07780029200280c1006;
assign testcases[239] = 76'h0778011a1002a0c1006;
assign testcases[240] = 76'h0788001a0001d0c0006;
assign testcases[241] = 76'h07780420701250c1006;
assign testcases[242] = 76'h07780119200240c1006;
assign testcases[243] = 76'h07780650a00451c1005;
assign testcases[244] = 76'h07780456600361c0005;
assign testcases[245] = 76'h19990991b0060473057;
assign testcases[246] = 76'h099a035190040283027;
assign testcases[247] = 76'h0cdc038d3001419104d;
assign testcases[248] = 76'h0ddd028d3000018104d;
assign testcases[249] = 76'h0ccc026d200170b001d;
assign testcases[250] = 76'h0bcc026d200251a101c;
assign testcases[251] = 76'h0aaa0b53700541c3007;
assign testcases[252] = 76'h18990652800551a3017;
assign testcases[253] = 76'h0778022910029190007;
assign testcases[254] = 76'h0788033920037181007;
assign testcases[255] = 76'h388907a2b0620706056;
assign testcases[256] = 76'h28790791b0320803026;
assign testcases[257] = 76'h887c0aa0c0400812026;
assign testcases[258] = 76'h28892ba0c0200803046;
assign testcases[259] = 76'h2879335290230704016;
assign testcases[260] = 76'h089924a880040322006;
assign testcases[261] = 76'h099905a880040323006;
assign testcases[262] = 76'h099908a880050431006;
assign testcases[263] = 76'h099905a880050421006;
assign testcases[264] = 76'h0889044930040421006;
assign testcases[265] = 76'h1bcb03aa70040245007;
assign testcases[266] = 76'h0899055280030273065;
assign testcases[267] = 76'h0899044180030273025;
assign testcases[268] = 76'h0999025a30020181026;
assign testcases[269] = 76'h0899024280030181026;
assign testcases[270] = 76'h0888014840110256075;
assign testcases[271] = 76'h0889034930000253055;
assign testcases[272] = 76'h07882a3180042261015;
assign testcases[273] = 76'h0788033270050240005;
assign testcases[274] = 76'h0788043170026170005;
assign testcases[275] = 76'h0788023270040251015;
assign testcases[276] = 76'h0788043170034260005;
assign testcases[277] = 76'h0888043a20032193015;
assign testcases[278] = 76'h0788012a20021181005;
assign testcases[279] = 76'h17883670a0231388034;
assign testcases[280] = 76'h08880991b0032294024;
assign testcases[281] = 76'h17780570a0220564024;
assign testcases[282] = 76'h199a046760250272018;
assign testcases[283] = 76'h0999035a30060270008;
assign testcases[284] = 76'h099a057950020271027;
assign testcases[285] = 76'h0bbb035c200260c000b;
assign testcases[286] = 76'h0bbb034c200290d000b;
assign testcases[287] = 76'h0aab036b300311a000b;
assign testcases[288] = 76'h0aaa036b300301a000b;
assign testcases[289] = 76'h0bbb024e1001a0d000b;
assign testcases[290] = 76'h0abb025c200340b000b;
assign testcases[291] = 76'h0aaa0b43700491a000b;
assign testcases[292] = 76'h0aaa0b71a006128000b;
assign testcases[293] = 76'h0aab0951900561a000b;
assign testcases[294] = 76'h0abb0594a00471c000c;
assign testcases[295] = 76'h0abb0494a004a1d000c;
assign testcases[296] = 76'h0bbb004d1001e0d010c;
assign testcases[297] = 76'h0bbb014e0001f0d000c;
assign testcases[298] = 76'h0bbb014d1001c0c000c;
assign testcases[299] = 76'h0bbb014d1001a0d000c;
assign testcases[300] = 76'h0aab014d100290d000b;
assign testcases[301] = 76'h0aab024d1001b0e000b;
assign testcases[302] = 76'h0aab014c100240d000b;
assign testcases[303] = 76'h0aab039c500270d010c;
assign testcases[304] = 76'h0abb014c200280e000c;
assign testcases[305] = 76'h0aab029c500350d010c;
assign testcases[306] = 76'h0abb014c200280e000c;
assign testcases[307] = 76'h0999013b100260a0008;
assign testcases[308] = 76'h0aab02337003c0d000a;
assign testcases[309] = 76'h0aab013d1001d0e000a;
assign testcases[310] = 76'h0bbc055a400381c000c;
assign testcases[311] = 76'h0bbb024c1001a0e000c;
assign testcases[312] = 76'h0bbc046c300361b000c;
assign testcases[313] = 76'h0abb045a300270d000c;
assign testcases[314] = 76'h0abb044a2002b0e000c;
assign testcases[315] = 76'h0abb015d200240c000c;
assign testcases[316] = 76'h0bbb045c2002a0d010d;
assign testcases[317] = 76'h0bbb014e0001f0e000d;
assign testcases[318] = 76'h0bbb045c2002a0d010b;
assign testcases[319] = 76'h0bbb014e0001f0e000d;
assign testcases[320] = 76'h0bbb005d100230d000d;
assign testcases[321] = 76'h0bbb034b200280d000d;
assign testcases[322] = 76'h0aaa075280057290009;
assign testcases[323] = 76'h0aaa03638002c1b0009;
assign testcases[324] = 76'h0aaa03638002c1b0009;
assign testcases[325] = 76'h1aab09a2c0052290119;
assign testcases[326] = 76'h0aab03437003b0e000b;
assign testcases[327] = 76'h0abb024d1001c0d000b;
assign testcases[328] = 76'h0abb014d1001e0f000c;
assign testcases[329] = 76'h0aaa014d100170e000c;
assign testcases[330] = 76'h0aab014d1001a0e000c;
assign testcases[331] = 76'h0aab014d1001a0e000c;
assign testcases[332] = 76'h0aaa004d100240e000c;
assign testcases[333] = 76'h0aab03437003b0e000b;
assign testcases[334] = 76'h0aab02437002e0e000b;
assign testcases[335] = 76'h0aab014d1001c0f000c;
assign testcases[336] = 76'h0aaa0243700321b0109;
assign testcases[337] = 76'h0aab014c200320b0009;
assign testcases[338] = 76'h0aab014c200320b0009;
assign testcases[339] = 76'h0999012c0001f0d0008;
assign testcases[340] = 76'h0999012c0001f0d0008;
assign testcases[341] = 76'h0999012c0001e0d0008;
assign testcases[342] = 76'h0999012c0001f0d0008;
assign testcases[343] = 76'h09aa0532700380d000a;
assign testcases[344] = 76'h0aaa213b100270e000a;
assign testcases[345] = 76'h09aa013c1001a0e000a;
assign testcases[346] = 76'h09aa013c1001a0e000a;
assign testcases[347] = 76'h09aa213b100220e000a;
assign testcases[348] = 76'h0aaa013c1001b0e100a;
assign testcases[349] = 76'h0aaa013d100290e100a;
assign testcases[350] = 76'h0aaa013d100190d000a;
assign testcases[351] = 76'h0aaa013d0001e0e000a;
assign testcases[352] = 76'h09aa013d0001f0e000a;
assign testcases[353] = 76'h0aaa024c200340c000a;
assign testcases[354] = 76'h09aa013b201240c000a;
assign testcases[355] = 76'h19aa28a2b03432a000a;
assign testcases[356] = 76'h0aaa0447500331a0007;
assign testcases[357] = 76'h099a075180050270017;
assign testcases[358] = 76'h099a0443700421a2008;
assign testcases[359] = 76'h09aa024370040191008;
assign testcases[360] = 76'h099a023c100240b1008;
assign testcases[361] = 76'h099a013c100250c1008;
assign testcases[362] = 76'h099a043a2002c0c1009;
assign testcases[363] = 76'h099a013c1001e0c1009;
assign testcases[364] = 76'h099a013c1001f0c1009;
assign testcases[365] = 76'h099a0439300341a1009;
assign testcases[366] = 76'h099a013c0001b0b1009;
assign testcases[367] = 76'h099a033a2002c0b1009;
assign testcases[368] = 76'h0999013b100211a1008;
assign testcases[369] = 76'h0aab025a302250b1009;
assign testcases[370] = 76'h0aab014b200240c0009;
assign testcases[371] = 76'h0aab044840130191009;
assign testcases[372] = 76'h1aab0458501261a1009;
assign testcases[373] = 76'h0aab024a301240c0009;
assign testcases[374] = 76'h0aab0348401321a1009;
assign testcases[375] = 76'h0bbc035a301270a100a;
assign testcases[376] = 76'h1bbc0c81b012529114a;
assign testcases[377] = 76'h0bbc0671a001027003a;
assign testcases[378] = 76'h0bbc035a301271a101a;
assign testcases[379] = 76'h0bbc047a4012319101a;
assign testcases[380] = 76'h0bbb0671a011028103a;
assign testcases[381] = 76'h4ab924b2c0010262177;
assign testcases[382] = 76'h4aca24b2c0010351167;
assign testcases[383] = 76'h29ba019b60010170127;
assign testcases[384] = 76'h0999014b20020180018;
assign testcases[385] = 76'h9acf3aa2c0160352167;
assign testcases[386] = 76'h6edf23a790000351137;
assign testcases[387] = 76'h8bcf07a690030251027;
assign testcases[388] = 76'h1998335190040260017;
assign testcases[389] = 76'hbabf66a1c0040351127;
assign testcases[390] = 76'h3aba54a1c0030351147;
assign testcases[391] = 76'h0abb245a300351a100b;
assign testcases[392] = 76'h0aab014d100290c000b;
assign testcases[393] = 76'h0bbb2493a004027100b;
assign testcases[394] = 76'h0abb2493a004219100b;
assign testcases[395] = 76'h0abb245a300361b100b;
assign testcases[396] = 76'h0abb2593a004218100b;
assign testcases[397] = 76'h0ccc016d200240b000c;
assign testcases[398] = 76'h0ccc006e100240b000c;
assign testcases[399] = 76'h1ccc07a0d024237001d;
assign testcases[400] = 76'h0cdd006f1001b19000d;
assign testcases[401] = 76'h0ccc04a2c012327000d;
assign testcases[402] = 76'h0ccc006f0001c18000d;
assign testcases[403] = 76'h0ccc006f0001c17000d;
assign testcases[404] = 76'h2bbc07b0d03282d000d;
assign testcases[405] = 76'h3bbc09b0d03183c000d;
assign testcases[406] = 76'h0bcc015e100290e000d;
assign testcases[407] = 76'h0bcc015e100250e000d;
assign testcases[408] = 76'h0bcc015b301280e000d;
assign testcases[409] = 76'h0bcc005e100290e000d;
assign testcases[410] = 76'h0abb0144700230c100c;
assign testcases[411] = 76'h0aba004d101230d100c;
assign testcases[412] = 76'h0bbb004e100220a000c;
assign testcases[413] = 76'h0bbb0144700320b000c;
assign testcases[414] = 76'h09aa0393a00311a1019;
assign testcases[415] = 76'h09a9024c20020190009;
assign testcases[416] = 76'h0aaa016c300211b0019;
assign testcases[417] = 76'h0aaa03bc600280c1019;
assign testcases[418] = 76'h0aaa014c1001c0d0009;
assign testcases[419] = 76'h0aab04bb700221b1019;
assign testcases[420] = 76'h0aaa03bc600180c0019;
assign testcases[421] = 76'h0abb045a300421b300b;
assign testcases[422] = 76'h0abb2653700451b100b;
assign testcases[423] = 76'h0aaa224c200301b100b;
assign testcases[424] = 76'h0abb245c200411b100b;
assign testcases[425] = 76'h0cdd226d2003119100f;
assign testcases[426] = 76'h0cdd03a88006119300f;
assign testcases[427] = 76'h1999245380020362094;
assign testcases[428] = 76'h089926b890020361054;
assign testcases[429] = 76'h089927b3c0020361064;
assign testcases[430] = 76'h0999264380020261074;
assign testcases[431] = 76'h099a045750040260066;
assign testcases[432] = 76'h189823a3b0040350056;
assign testcases[433] = 76'h099a035a30020270036;
assign testcases[434] = 76'h3cbc57b0d07343b500d;
assign testcases[435] = 76'h2bbc0770b02132a200d;
assign testcases[436] = 76'h2cbc3ab0d04152b300d;
assign testcases[437] = 76'h2bbc27b0d04333a400d;
assign testcases[438] = 76'h3cbcdbb0d04936a400d;
assign testcases[439] = 76'h4bbcbab0d047169300d;
assign testcases[440] = 76'h1aab5b60a025239101b;
assign testcases[441] = 76'h1aab5d60a023239101b;
assign testcases[442] = 76'h1bbb0361a01311a000b;
assign testcases[443] = 76'h0bbb005d100210a000b;
assign testcases[444] = 76'h0bbb016d200211a000b;
assign testcases[445] = 76'h0aaa014d100270c000b;
assign testcases[446] = 76'h0aaa014d100270c000b;
assign testcases[447] = 76'h0aaa014d100270c000b;
assign testcases[448] = 76'h0aaa0463800221a0039;
assign testcases[449] = 76'h09aa0463800331a0019;
assign testcases[450] = 76'h09aa0449300331a0009;
assign testcases[451] = 76'h0aaa0463800111a0039;
assign testcases[452] = 76'h19990991b0060473066;
assign testcases[453] = 76'h099a013b20033191008;
assign testcases[454] = 76'h099a023b200331a1008;
assign testcases[455] = 76'h099a023b20032191008;
assign testcases[456] = 76'h1999025090160553147;
assign testcases[457] = 76'h1bbc2793a005046104a;
assign testcases[458] = 76'h0bbc01739005027002a;
assign testcases[459] = 76'h0aba03639003117102a;
assign testcases[460] = 76'h07780238300220b1024;
assign testcases[461] = 76'h06780229100240c0004;
assign testcases[462] = 76'h0788013830030191024;
assign testcases[463] = 76'h18872e71a0041381044;
assign testcases[464] = 76'h1787066380031191014;
assign testcases[465] = 76'h0abb04b4b01341e100b;
assign testcases[466] = 76'h0aab027c300250f100b;
assign testcases[467] = 76'h0aab027c300250f100b;
assign testcases[468] = 76'h0aab027c300260f100b;
assign testcases[469] = 76'h0bcc026c300250f000d;
assign testcases[470] = 76'h0bbc025c200250f000d;
assign testcases[471] = 76'h0bcc005e100270f000d;
assign testcases[472] = 76'h0bbc027c400230f100d;
assign testcases[473] = 76'h0bcb017b400340f000d;
assign testcases[474] = 76'h0bbb005d200260f000d;
assign testcases[475] = 76'h0bbb005d100270f000d;
assign testcases[476] = 76'h0abb2153801311b100c;
assign testcases[477] = 76'h0bbb015c200220c000c;
assign testcases[478] = 76'h0abb2159401211a100c;
assign testcases[479] = 76'h0bbb2159401201a000c;
assign testcases[480] = 76'h0aaa08b4b00461a100a;
assign testcases[481] = 76'h0aaa0455700271b000a;
assign testcases[482] = 76'h0abb269b5003119001a;
assign testcases[483] = 76'h1abc2571b003129001a;
assign testcases[484] = 76'h0aab2954700531a100b;
assign testcases[485] = 76'h0aab024d100230b000b;
assign testcases[486] = 76'h28a90582a0120250066;
assign testcases[487] = 76'h29a90582b0010250046;
assign testcases[488] = 76'h2899047480120340026;
assign testcases[489] = 76'h29a90582a0010250066;
assign testcases[490] = 76'h4cbd0971b0040551284;
assign testcases[491] = 76'h5cbd08a0d0030640164;
assign testcases[492] = 76'h3cbd0ca0c0000451264;
assign testcases[493] = 76'h2ccd0580b0030451244;
assign testcases[494] = 76'h2aa92c72a0020551176;
assign testcases[495] = 76'h39a92572a0020361146;
assign testcases[496] = 76'h2bbc0970b00305413a7;
assign testcases[497] = 76'h1bbc0780c0010451267;
assign testcases[498] = 76'h1cbc0b70b0040640387;
assign testcases[499] = 76'h2bbc0980c0020451277;
assign testcases[500] = 76'h2bab2a70b00208411a7;
assign testcases[501] = 76'h1bab2990c0020741077;
assign testcases[502] = 76'h2bbc0571a0060453067;
assign testcases[503] = 76'h2bbc0470a0050453047;
assign testcases[504] = 76'h19a90681b0040262047;
assign testcases[505] = 76'h19a90781b0040262027;
assign testcases[506] = 76'h0ded00af3002018106f;
assign testcases[507] = 76'h0ded01af3002018104f;
assign testcases[508] = 76'h0ded01af3002018105f;
assign testcases[509] = 76'h1ded02af3001018103f;
assign testcases[510] = 76'h0ddd339b6002018204e;
assign testcases[511] = 76'h1ded229e4001017104e;
assign testcases[512] = 76'h0cdd017d3003019101e;
assign testcases[513] = 76'h0cdd218f2002019001e;
assign testcases[514] = 76'h1aa9245380020274167;
assign testcases[515] = 76'h19a9035380020172127;
assign testcases[516] = 76'h19a9038490010262037;
assign testcases[517] = 76'h1aac0383a0010272147;
assign testcases[518] = 76'h189908a2b0030363146;
assign testcases[519] = 76'h189908a0d0020362136;
assign testcases[520] = 76'h0889034280041261016;
assign testcases[521] = 76'h0889213a20031260006;
assign testcases[522] = 76'h1fff04af4004026116f;
assign testcases[523] = 76'h1fff02af4000016114f;
assign testcases[524] = 76'h1fff01af3000026114f;
assign testcases[525] = 76'h1fff02af4001026003f;
assign testcases[526] = 76'h3edf0bb0d01104512bb;
assign testcases[527] = 76'h1fef079b5000036116b;
assign testcases[528] = 76'h1fff02997000026114b;
assign testcases[529] = 76'h2cce09b1d000054014b;
assign testcases[530] = 76'h3ccd09b0d011074014b;
assign testcases[531] = 76'h1fff04a3b000036116b;
assign testcases[532] = 76'h0aaa0763800441a0029;
assign testcases[533] = 76'h0aaa0363800441a0009;
assign testcases[534] = 76'h0aaa0363800261b0009;
assign testcases[535] = 76'h0aaa277490053290019;
assign testcases[536] = 76'h0aaa047490024190019;
assign testcases[537] = 76'h0aab0463800551b000b;
assign testcases[538] = 76'h0aab0463800451c000b;
assign testcases[539] = 76'h0aaa0461a00341b000b;
assign testcases[540] = 76'h0ccc04648003018104c;
assign testcases[541] = 76'h0ccc006e2002019001c;
assign testcases[542] = 76'h0abb06619005019101a;
assign testcases[543] = 76'h0aba04537005019100a;
assign testcases[544] = 76'h0abb044b201250c000c;
assign testcases[545] = 76'h0abb014d100270c100c;
assign testcases[546] = 76'h0aab044b300340b000c;
assign testcases[547] = 76'h0abb0447501251a2109;
assign testcases[548] = 76'h0aab014c200331a300a;
assign testcases[549] = 76'h0aab014c100240a100a;
assign testcases[550] = 76'h0aab014b200241a200a;
assign testcases[551] = 76'h4bbb54b0d0090d55079;
assign testcases[552] = 76'h4cdb3ab0d0020b52079;
assign testcases[553] = 76'h3aab2970b0490b5702a;
assign testcases[554] = 76'h2a9a2880b047095300a;
assign testcases[555] = 76'h3bbb27b0d00b0c6302a;
assign testcases[556] = 76'h1aaa0480b037086401a;
assign testcases[557] = 76'h299935a0d0290662027;
assign testcases[558] = 76'h289936a0d0230552027;
assign testcases[559] = 76'h389827a0d0240651017;
assign testcases[560] = 76'h1778244180210450007;
assign testcases[561] = 76'h288928a1c0350658017;
assign testcases[562] = 76'h17792760a0340474007;
assign testcases[563] = 76'h479809a0c0250745017;
assign testcases[564] = 76'h589828a1c0160833017;
assign testcases[565] = 76'h19992880b0430674057;
assign testcases[566] = 76'h18892ab0d0410572037;
assign testcases[567] = 76'h199907a0c0221483037;
assign testcases[568] = 76'h18893bb0d0410563037;
assign testcases[569] = 76'h489935a0d0650856057;
assign testcases[570] = 76'h18890580b0460663017;
assign testcases[571] = 76'h59a926b0d0360853047;
assign testcases[572] = 76'h59a936a0d0460854047;
assign testcases[573] = 76'h69b926b0d0180953037;
assign testcases[574] = 76'h8dc936b0d0150b51037;
assign testcases[575] = 76'h18792480b0450663007;
assign testcases[576] = 76'h18890680b0450663017;
assign testcases[577] = 76'h09aa0481b01501c0029;
assign testcases[578] = 76'h2798057860030263024;
assign testcases[579] = 76'h0778022920040171004;
assign testcases[580] = 76'h0888012920030251014;
assign testcases[581] = 76'h1788047860030263024;
assign testcases[582] = 76'h2798047960030261014;
assign testcases[583] = 76'h2798067960030263024;
assign testcases[584] = 76'h16770971a0140262014;
assign testcases[585] = 76'h0667033830130271004;
assign testcases[586] = 76'h0678012820040261004;
assign testcases[587] = 76'h27870572a0040353124;
assign testcases[588] = 76'h0677056850050361004;
assign testcases[589] = 76'h0677046850050361004;
assign testcases[590] = 76'h38980692b0030453124;
assign testcases[591] = 76'h49ad247770050352014;
assign testcases[592] = 76'h49ad067480010352024;
assign testcases[593] = 76'h3797047480040352024;
assign testcases[594] = 76'h0bcb027d300311e301c;
assign testcases[595] = 76'h0bbb015d200310e300c;
assign testcases[596] = 76'h0bbb005e100310f200c;
assign testcases[597] = 76'h0bbb017d300311e200c;
assign testcases[598] = 76'h0bbb017d300311e300c;
assign testcases[599] = 76'h0bbb017d300301d100c;
assign testcases[600] = 76'h0bcc0475801301d104b;
assign testcases[601] = 76'h0bcc028b500401e101b;
assign testcases[602] = 76'h0bcc0375801101d104b;
assign testcases[603] = 76'h0ccc0385901201d104b;
assign testcases[604] = 76'h0bbb0473900302c002b;
assign testcases[605] = 76'h1ccc02aa700301d206c;
assign testcases[606] = 76'h1ccc01aa600301c102c;
assign testcases[607] = 76'h1cdc02aa700301d204c;
assign testcases[608] = 76'h1bbb24739006035204b;
assign testcases[609] = 76'h1bbb2271a004035103b;
assign testcases[610] = 76'h1bbb2571a008045101b;
assign testcases[611] = 76'h1bbb24739007044103b;
assign testcases[612] = 76'h0bbb28a1c003036101b;
assign testcases[613] = 76'h1bcc0680b009046107c;
assign testcases[614] = 76'h1bbc0470b008046105c;
assign testcases[615] = 76'h1ccc0780c008046104c;
assign testcases[616] = 76'h1ddc0393a000026118c;
assign testcases[617] = 76'h1aaa0150900c164100b;
assign testcases[618] = 76'h0aab02418003226000b;
assign testcases[619] = 76'h1bcb0480c003027306b;
assign testcases[620] = 76'h1ccc0490c001027206b;
assign testcases[621] = 76'h0abb026d2003117100b;
assign testcases[622] = 76'h2a9a045190090753168;
assign testcases[623] = 76'h199a0361a0060561048;
assign testcases[624] = 76'h19990260a0090672157;
assign testcases[625] = 76'h19a90260a0090572147;
assign testcases[626] = 76'h2aaa0960a0150550038;
assign testcases[627] = 76'h17780891c0162371024;
assign testcases[628] = 76'h0778002a20025181004;
assign testcases[629] = 76'h2bbb0471a03006730a8;
assign testcases[630] = 76'h2bbd0470b0000582098;
assign testcases[631] = 76'h0bbc0893a007228000b;
assign testcases[632] = 76'h0bbc24648004217000b;
assign testcases[633] = 76'h0bcc015e100211b000b;
assign testcases[634] = 76'h0bbb07b4b014128002b;
assign testcases[635] = 76'h0bbb0274900311a000b;
assign testcases[636] = 76'h0bbb03685003019000b;
assign testcases[637] = 76'h0abb05849004037002b;
assign testcases[638] = 76'h0aab0693a0040270039;
assign testcases[639] = 76'h0aab0493a0040260029;
assign testcases[640] = 76'h0aab045370050260009;
assign testcases[641] = 76'h0aab035380060260009;
assign testcases[642] = 76'h1aab8490c0060560069;
assign testcases[643] = 76'h0abb0bb0d0020370049;
assign testcases[644] = 76'h077803292002d0d1005;
assign testcases[645] = 76'h0778011a1001f0e0005;
assign testcases[646] = 76'h07780425400301a1005;
assign testcases[647] = 76'h077803254002b0d1005;
assign testcases[648] = 76'h077803254002a0d1005;
assign testcases[649] = 76'h077801172002c0c0005;
assign testcases[650] = 76'h0778021a1001f0d0005;
assign testcases[651] = 76'h0778021a1001f0d0005;
assign testcases[652] = 76'h07780017300290c0005;
assign testcases[653] = 76'h077802191001c0c0005;
assign testcases[654] = 76'h077801191001e0d0005;
assign testcases[655] = 76'h0899065280032324027;
assign testcases[656] = 76'h09990882a0031323027;
assign testcases[657] = 76'h0899024a30022323017;
assign testcases[658] = 76'h0999015a30022232017;
assign testcases[659] = 76'h0899014a30022322017;
assign testcases[660] = 76'h0899024a30022322017;
assign testcases[661] = 76'h624439a0d4500e21007;
assign testcases[662] = 76'h498a28a1c81323a3009;
assign testcases[663] = 76'h498a2aa1c81323a3009;
assign testcases[664] = 76'h498a2993a40212a1009;
assign testcases[665] = 76'h398a2b93a40322a2009;
assign testcases[666] = 76'h0aaa014a200321b1009;
assign testcases[667] = 76'h0aaa034c200220b1009;
assign testcases[668] = 76'h399a37a1c41232a2009;
assign testcases[669] = 76'h3aab3b91b033129101a;
assign testcases[670] = 76'h4a9b37a1c033229101a;
assign testcases[671] = 76'h1aac25585013017000a;
assign testcases[672] = 76'h0bbb015b300221b101a;
assign testcases[673] = 76'h2ddf0490c00103a109a;
assign testcases[674] = 76'h2edf0490c00303a106a;
assign testcases[675] = 76'h2ddb0390c000039006a;
assign testcases[676] = 76'h2edf018a500002a004a;
assign testcases[677] = 76'h2ddf0390c000039006a;
assign testcases[678] = 76'h2edf0492b00102a004a;
assign testcases[679] = 76'h0aab07619008028301b;
assign testcases[680] = 76'h0abb037a4003019101b;
assign testcases[681] = 76'h1abb3882a00d065302a;
assign testcases[682] = 76'h602238b1d8200651508;
assign testcases[683] = 76'h50222461a8100551408;
assign testcases[684] = 76'h199a015660250336528;
assign testcases[685] = 76'h199a025380240334428;
assign testcases[686] = 76'h0999013930050341008;
assign testcases[687] = 76'h199a025660240333328;
assign testcases[688] = 76'h199a025380130333428;
assign testcases[689] = 76'h598a067294450523e38;
assign testcases[690] = 76'h3677047294170611508;
assign testcases[691] = 76'h299a267390240431828;
assign testcases[692] = 76'h498a0580b0340432838;
assign testcases[693] = 76'h28892681a4430444f38;
assign testcases[694] = 76'h1999065380220352928;
assign testcases[695] = 76'h2879045194320433918;
assign testcases[696] = 76'h1999045380130342828;
assign testcases[697] = 76'h67690c61a8430443d17;
assign testcases[698] = 76'h94422981b4210551607;
assign testcases[699] = 76'h28890ea1c4430432917;
assign testcases[700] = 76'h87590c91cc320542907;
assign testcases[701] = 76'h38790a91b41404a1507;
assign testcases[702] = 76'h37860337440200f0307;
assign testcases[703] = 76'h27760337440200f0307;
assign testcases[704] = 76'h16760128240000f0207;
assign testcases[705] = 76'h089927b3b003a1a6008;
assign testcases[706] = 76'h0899012b1001e0b4008;
assign testcases[707] = 76'h0899023a20031196017;
assign testcases[708] = 76'h0899013b20022193007;
assign testcases[709] = 76'h0889023a20025194006;
assign testcases[710] = 76'h0889023a20027191006;
assign testcases[711] = 76'h18892770b0280463026;
assign testcases[712] = 76'h1889044090070462026;
assign testcases[713] = 76'h1889075090061371024;
assign testcases[714] = 76'h09a9025a40033195048;
assign testcases[715] = 76'h0aaa025a40030193038;
assign testcases[716] = 76'h0899025a300241a3018;
assign testcases[717] = 76'h0899023a200270b1008;
assign testcases[718] = 76'h099a225a30040181018;
assign testcases[719] = 76'h0889013a200290b3007;
assign testcases[720] = 76'h0889012b0001d0b1007;
assign testcases[721] = 76'h0abb025c200280b010b;
assign testcases[722] = 76'h0abb015e100290c000b;
assign testcases[723] = 76'h0abb045a4004119010b;
assign testcases[724] = 76'h09aa045a30020192147;
assign testcases[725] = 76'h09aa035a30020192027;
assign testcases[726] = 76'h09aa035750030191007;
assign testcases[727] = 76'h19a9005a30010191027;
assign testcases[728] = 76'h0788024180021183024;
assign testcases[729] = 76'h1788024180021182024;
assign testcases[730] = 76'h0778012a10031191004;
assign testcases[731] = 76'h2aac025a40030171024;
assign testcases[732] = 76'h0788034a30021182014;
assign testcases[733] = 76'h1bbb289a60030366165;
assign testcases[734] = 76'h1aab0594a0020271147;
assign testcases[735] = 76'h1bbb299a60020363167;
assign testcases[736] = 76'h1bbb289a60030364147;
assign testcases[737] = 76'h1888063180070463065;
assign testcases[738] = 76'h1889253080050361045;
assign testcases[739] = 76'h1778246190081561044;
assign testcases[740] = 76'h1889046190060460044;
assign testcases[741] = 76'h0abb02629002119102a;
assign testcases[742] = 76'h0abb015d100210a101a;
assign testcases[743] = 76'h398a3790c0b1073301b;
assign testcases[744] = 76'h56655c80b0500a0100b;
assign testcases[745] = 76'h498a2ba0d091082301b;
assign testcases[746] = 76'h299a07a0d081064301b;
assign testcases[747] = 76'h398a06a0d081073301b;
assign testcases[748] = 76'h0999023b100270e0008;
assign testcases[749] = 76'h0999023c100290f0008;
assign testcases[750] = 76'h0999013c1001b0f0008;
assign testcases[751] = 76'h0999023b100270e0008;
assign testcases[752] = 76'h0899048b50026190017;
assign testcases[753] = 76'h0899023b10026190007;
assign testcases[754] = 76'h0899013b200260a0007;
assign testcases[755] = 76'h0899023b200270a0007;
assign testcases[756] = 76'h0889033080071270007;
assign testcases[757] = 76'h0889012260042280007;
assign testcases[758] = 76'h08992692b00301a0027;
assign testcases[759] = 76'h0899003b200300c0007;
assign testcases[760] = 76'h09aa0489600210a0027;
assign testcases[761] = 76'h099a024a200210a0027;
assign testcases[762] = 76'h099a004b200220c0007;
assign testcases[763] = 76'h09990f92a00642a0027;
assign testcases[764] = 76'h0aaa0243700380c000a;
assign testcases[765] = 76'h0aaa013c1001b0e000a;
assign testcases[766] = 76'h0aab014c100250a000a;
assign testcases[767] = 76'h099a02327001c0c0009;
assign testcases[768] = 76'h099a013c1001d0c0009;
assign testcases[769] = 76'h0999012c0000f0f0008;
assign testcases[770] = 76'h0999012c0000f0f0008;
assign testcases[771] = 76'h088905282011f0e0007;
assign testcases[772] = 76'h08890568501170d0007;
assign testcases[773] = 76'h0889012b0001f0e0007;
assign testcases[774] = 76'h088905685011c0d0007;
assign testcases[775] = 76'h09aa025b200270e1009;
assign testcases[776] = 76'h09aa024b200260d1009;
assign testcases[777] = 76'h09aa024b200260d1009;
assign testcases[778] = 76'h09aa024b200250d1009;
assign testcases[779] = 76'h0899013b200260d0007;
assign testcases[780] = 76'h0889013b200270d0007;
assign testcases[781] = 76'h0999023b100260e0007;
assign testcases[782] = 76'h0889013b200280d0007;
assign testcases[783] = 76'h0999049b500340c0008;
assign testcases[784] = 76'h0999023a300340d0008;
assign testcases[785] = 76'h0778052170041190013;
assign testcases[786] = 76'h0778042170042180003;
assign testcases[787] = 76'h0889062080050190025;
assign testcases[788] = 76'h0888062270051190025;
assign testcases[789] = 76'h0888044560020190015;
assign testcases[790] = 76'h0889062170051280015;
assign testcases[791] = 76'h0889062170051280015;
assign testcases[792] = 76'h0bbb04666053619c01c;
assign testcases[793] = 76'h1bbc03666053619901c;
assign testcases[794] = 76'h1bbc03657053628801c;
assign testcases[795] = 76'h0bbb025d100250b400c;
assign testcases[796] = 76'h0bbb015d100260c300c;
assign testcases[797] = 76'h0bbb015d100270b300c;
assign testcases[798] = 76'h0bbb015d100270b300c;
assign testcases[799] = 76'h0bbc035c200280b400c;
assign testcases[800] = 76'h0bbc005e1001a0c300c;
assign testcases[801] = 76'h0bbc046c201270b500c;
assign testcases[802] = 76'h0bbb016c200260b300c;
assign testcases[803] = 76'h2aab04657052343200c;
assign testcases[804] = 76'h1aab03657054243301c;
assign testcases[805] = 76'h0ccd036a4003518100c;
assign testcases[806] = 76'h0ccd226d2003619100c;
assign testcases[807] = 76'h0ccd226d2003619100c;
assign testcases[808] = 76'h1cbc22758052626402c;
assign testcases[809] = 76'h0ccc046a400290a100c;
assign testcases[810] = 76'h0ccc24666013819100c;
assign testcases[811] = 76'h1ccd32767032535302c;
assign testcases[812] = 76'h1ccd52767022626302c;
assign testcases[813] = 76'h2cbd21758042434302c;
assign testcases[814] = 76'h2bbb04748022033101c;
assign testcases[815] = 76'h1bbb04647022333100c;
assign testcases[816] = 76'h1bbb04647022333101c;
assign testcases[817] = 76'h0ccd026b3003a0a100e;
assign testcases[818] = 76'h0ccd026b300391a100e;
assign testcases[819] = 76'h0ccd236c3002b0a200e;
assign testcases[820] = 76'h0ccd236c3002a0a100e;
assign testcases[821] = 76'h0ccd016f1001c0b200e;
assign testcases[822] = 76'h0ccd016f1001b0a200e;
assign testcases[823] = 76'h0ccd046c2002c0a200e;
assign testcases[824] = 76'h0ccd046b3002d0a100e;
assign testcases[825] = 76'h0ccc005d2002a0b300e;
assign testcases[826] = 76'h0ccc5469501281a300e;
assign testcases[827] = 76'h0ccc54676012819200e;
assign testcases[828] = 76'h0ccd236b3003b1a200e;
assign testcases[829] = 76'h0ccc33695012a1a300e;
assign testcases[830] = 76'h0ccc5469501291a300e;
assign testcases[831] = 76'h0ccc54575011b1a100e;
assign testcases[832] = 76'h0ccc33575012719300e;
assign testcases[833] = 76'h0ccd046b300381a100e;
assign testcases[834] = 76'h3aac267390510522047;
assign testcases[835] = 76'h298a2571a0510711027;
assign testcases[836] = 76'h2a9b227480440621017;
assign testcases[837] = 76'h3aac227480420531047;
assign testcases[838] = 76'h09aa03493002a173009;
assign testcases[839] = 76'h09aa03493002b173009;
assign testcases[840] = 76'h09aa044930029171009;
assign testcases[841] = 76'h0aaa034930028161009;
assign testcases[842] = 76'h0aaa024930028163009;
assign testcases[843] = 76'h0aaa014c1002b172009;
assign testcases[844] = 76'h0aaa014c10029172009;
assign testcases[845] = 76'h0aaa044840032162019;
assign testcases[846] = 76'h0aaa044840032163019;
assign testcases[847] = 76'h0aaa044840031163019;
assign testcases[848] = 76'h0aaa045840031163019;
assign testcases[849] = 76'h0aaa045840031163019;
assign testcases[850] = 76'h0aaa005c20032172019;
assign testcases[851] = 76'h0abb005c20022173019;
assign testcases[852] = 76'h0aaa024c20032161009;
assign testcases[853] = 76'h09aa024c20027161009;
assign testcases[854] = 76'h0aaa013c1002a171009;
assign testcases[855] = 76'h0aab015c2003417200b;
assign testcases[856] = 76'h0aab015c2003117100b;
assign testcases[857] = 76'h0abb015b3004017300b;
assign testcases[858] = 76'h0abb005b3004016300b;
assign testcases[859] = 76'h0bbb005b3004026100b;
assign testcases[860] = 76'h0bbb015b3004026201b;
assign testcases[861] = 76'h0bbb015c2002517201b;
assign testcases[862] = 76'h0abb04638004225201b;
assign testcases[863] = 76'h0abb035c2002717301b;
assign testcases[864] = 76'h0bbb005c2003317101b;
assign testcases[865] = 76'h0bbb015b3004026101b;
assign testcases[866] = 76'h0bbb015d1002518100b;
assign testcases[867] = 76'h0abb035c2002717301b;
assign testcases[868] = 76'h0abb045a3002717301b;
assign testcases[869] = 76'h0aaa025a30014164059;
assign testcases[870] = 76'h0aaa225a30014163049;
assign testcases[871] = 76'h0aaa025a30013162029;
assign testcases[872] = 76'h0aaa035a30014163029;
assign testcases[873] = 76'h0aaa015c20013172019;
assign testcases[874] = 76'h0aaa024b20022172019;
assign testcases[875] = 76'h0aaa034a30031163019;
assign testcases[876] = 76'h0aaa034a30031163019;
assign testcases[877] = 76'h09aa024a30031163019;
assign testcases[878] = 76'h09aa014840041263019;
assign testcases[879] = 76'h09aa024a30040253019;
assign testcases[880] = 76'h09aa024840040252019;
assign testcases[881] = 76'h09aa034930040263009;
assign testcases[882] = 76'h09aa024b20030253019;
assign testcases[883] = 76'h09aa035b30032253019;
assign testcases[884] = 76'h09aa045b30025162019;
assign testcases[885] = 76'h0aaa013c10028171009;
assign testcases[886] = 76'h0aaa024c10018173019;
assign testcases[887] = 76'h0aab014c10024183009;
assign testcases[888] = 76'h0aab014d10025192009;
assign testcases[889] = 76'h0aaa014d10018172019;
assign testcases[890] = 76'h0aaa014d10027173019;
assign testcases[891] = 76'h0aab014d10025183009;
assign testcases[892] = 76'h0aaa034c20027173019;
assign testcases[893] = 76'h0bbb015c2003116300b;
assign testcases[894] = 76'h0abb005c2003015400b;
assign testcases[895] = 76'h0bbb005c2004125400b;
assign testcases[896] = 76'h0bbb005b3003025501b;
assign testcases[897] = 76'h0bbb015b3004024300b;
assign testcases[898] = 76'h0bbb006b4004024301b;
assign testcases[899] = 76'h0bbb047a5004024201b;
assign testcases[900] = 76'h1bbb037a5006034201b;
assign testcases[901] = 76'h1bbb23777027033401b;
assign testcases[902] = 76'h1aab33777027042300b;
assign testcases[903] = 76'h0bbb25767017233500c;
assign testcases[904] = 76'h0abb04667026134500c;
assign testcases[905] = 76'h0aab03575031024300c;
assign testcases[906] = 76'h0bbb32685032024302c;
assign testcases[907] = 76'h0bbb22676022034302c;
assign testcases[908] = 76'h0bcc269a6002033606c;
assign testcases[909] = 76'h0ccc049b5003033302c;
assign testcases[910] = 76'h2aab27b0d055081001c;
assign testcases[911] = 76'h2bbc27748054053102c;
assign testcases[912] = 76'h0bcc047a5015033302c;
assign testcases[913] = 76'h0778011820032161005;
assign testcases[914] = 76'h0778021730030151005;
assign testcases[915] = 76'h0778233740030241015;
assign testcases[916] = 76'h1778213554010331015;
assign testcases[917] = 76'h1668343554021242005;
assign testcases[918] = 76'h1668021540122251005;
assign testcases[919] = 76'h0678011820032162005;
assign testcases[920] = 76'h0788022920032153005;
assign testcases[921] = 76'h0778022730231243005;
assign testcases[922] = 76'h1778223554030241015;
assign testcases[923] = 76'h0778223740030341015;
assign testcases[924] = 76'h1889024650220242025;
assign testcases[925] = 76'h1778035560231423015;
assign testcases[926] = 76'h0778043650141332005;
assign testcases[927] = 76'h1778025660320333015;
assign testcases[928] = 76'h1778033640330333015;
assign testcases[929] = 76'h1889024650220242025;
assign testcases[930] = 76'h0899234750030253025;
assign testcases[931] = 76'h0778012640340344005;
assign testcases[932] = 76'h0788012920040255005;
assign testcases[933] = 76'h1778035660231333015;
assign testcases[934] = 76'h188a034090250433016;
assign testcases[935] = 76'h089a233740130243016;
assign testcases[936] = 76'h0899013930040244006;
assign testcases[937] = 76'h0899013930050255006;
assign testcases[938] = 76'h0899013930050255006;
assign testcases[939] = 76'h199a546480226293009;
assign testcases[940] = 76'h0aaa014b2002b0c1009;
assign testcases[941] = 76'h09aa085b300381a3019;
assign testcases[942] = 76'h09aa065a40033193029;
assign testcases[943] = 76'h0bbb016a40031191029;
assign testcases[944] = 76'h37683560a8400531019;
assign testcases[945] = 76'h2bab5560a0213270029;
assign testcases[946] = 76'h1aab04547035134300b;
assign testcases[947] = 76'h1aab24547035034502b;
assign testcases[948] = 76'h0bbb34594004017103b;
assign testcases[949] = 76'h0bbb06585003016102b;
assign testcases[950] = 76'h0bbb24566006025402b;
assign testcases[951] = 76'h1abb02566008024100b;
assign testcases[952] = 76'h1aab045280320254069;
assign testcases[953] = 76'h199a025280430252039;
assign testcases[954] = 76'h199a035380440255009;
assign testcases[955] = 76'h199a066290460345009;
assign testcases[956] = 76'h1999046380640345009;
assign testcases[957] = 76'h1999244370530343009;
assign testcases[958] = 76'h199a044280350243009;
assign testcases[959] = 76'h398a065290670624008;
assign testcases[960] = 76'h487a065290660623008;
assign testcases[961] = 76'h199a065280391354008;
assign testcases[962] = 76'h298a054280941341018;
assign testcases[963] = 76'h198a044370651351008;
assign testcases[964] = 76'h299a244280460433038;
assign testcases[965] = 76'h299a344180350332018;
assign testcases[966] = 76'h199a384280170442028;
assign testcases[967] = 76'h199a384280160431028;
assign testcases[968] = 76'h199a285280190253008;
assign testcases[969] = 76'h099a375560091263008;
assign testcases[970] = 76'h099a023560162171008;
assign testcases[971] = 76'h4879266190911444007;
assign testcases[972] = 76'h587a266190711534007;
assign testcases[973] = 76'h4879235180611443007;
assign testcases[974] = 76'h2879043360411261007;
assign testcases[975] = 76'h598a256190522543007;
assign testcases[976] = 76'h299a054090412263017;
assign testcases[977] = 76'h399a064090322263007;
assign testcases[978] = 76'h598a0680b4710443027;
assign testcases[979] = 76'h5a8a2580b4300451027;
assign testcases[980] = 76'h4a9a044180410362027;
assign testcases[981] = 76'h1a9a024470210262027;
assign testcases[982] = 76'h0899004a30040243007;
assign testcases[983] = 76'h0899003a30040242007;
assign testcases[984] = 76'h099a004b20040241017;
assign testcases[985] = 76'h09aa015a40020333047;
assign testcases[986] = 76'h09aa025a40020333037;
assign testcases[987] = 76'h0aba077a40010334077;
assign testcases[988] = 76'h1aba077580010343057;
assign testcases[989] = 76'h0bbb037b40020323077;
assign testcases[990] = 76'h1aaa058580020331047;
assign testcases[991] = 76'h19aa046570020331047;
assign testcases[992] = 76'h0abb067a40030333067;
assign testcases[993] = 76'h0aba067580010333067;
assign testcases[994] = 76'h0899035750020231027;
assign testcases[995] = 76'h0899014b20020230017;
assign testcases[996] = 76'h1899046850140333047;
assign testcases[997] = 76'h19a9015a40040323047;
assign testcases[998] = 76'h19a9015940040332047;
assign testcases[999] = 76'h0aab046950000325087;


  
  localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
  wire [$clog2(CLASS_CNT)-1:0] prediction;

  // Instantiate module under test
 cardio_bnn1_bnnseq #() dut (
    .features(sample),
    .clk(clk),
    .rst(rst),
    .prediction(prediction)
  );
  
  always #halfPeriod clk <= ~clk;

  integer i;
  initial begin
    $write("["); //"
    for(i=0;i<TEST_CNT;i=i+1)
        runtestcase(i);
    $display("]");
    $finish;
  end

  localparam [$clog2(CLASS_CNT)-1:0] maxclass = CLASS_CNT-1;

  task runtestcase(input integer i); begin
    sample <= testcases[i];
    rst <= 1;
    clk <= 0;
    #period
    rst <= 0;
    #period
    #((FEAT_CNT+HIDDEN_CNT-1)*period)
    $write("%d, ",(prediction));
  end
  endtask

endmodule
