











module pendigits_tnn1_tnnzeq #(

parameter FEAT_CNT = 16,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 10,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnnzeq #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(640'b0100100000101010010010000000101001100001000010101001001000010001000100000000000010010010100000010100100100100101100010101111010001001101110000001011001010100101010110100000001110101001000010101111101100010000010010100101001010100000000110100000010000000110010000010011100010001011110100000110110110000010101000000000101010100100000110100001000000011010110000101011110010110000000011010100101000000000111010001111010010100001100000000100000101101000010000000000111011111000000100110001000001011000010010101100000010101100000001100001011000000001101000000010011000000000000110101110111110000101000100000101101010110010000000110101000001001001),
  .MASK(640'b1111100110101011111110101011111111110001100110111011001100010011101110011010010011011011100000111110100101101111101011111111010111001111111110101011101111111111111110110101111110111011001111111111111100011111010111111111111111111111100110101110111000010110111111110011101110011011110110111111110110011110111110101000101111111110101110110011101010011010111101111011111011111111010111011111101010000001111011011111111111101001100000001111111101101011110101110001111011111011101101111111100011111101111110101111000111111100100011101111111101000001111011101110011010100000100111111111111111011111111110100111111111110011010000111111110101101101),
  .NONZERO_CNT(640'h0b0d0a0808090b0c0c0e0d0c0d0e0c090d0b0c0a0d080d0d080e060d0a0d0c0b0a0a0b080f0d090c),
  .SPARSE_VALS2(208'b0111001101000010010001110110101010101100000001110111100101000001100011101000110111110011111010001010111010111000100010011010000011011010101010110100110011011100010101011001000111100100000000100010000010100101),  // Bits of not-zeroes
  .COL_INDICES(1664'h25201f1e191716151311100f0c070605040327252322201e1d1c1b1a191817151211100f0e0d0b080604241f1d1c1b191817150e0c0706040302002522201b191817161514131211100f0e0c0b0a080706050127231f1e1a1816110f0e0c0a0907020100272321201f1e1d1c1b1a1716151413110f0e0d0b0a0503021f1e1d1c171615130f0e0c0a090806050403020100271e1c191714130f0e0d0c0b0807060504030201002321201c1a17161312110f0e0c0a0908070605010027201d1b1817161312110e0c0b0a08070504030201), // Column of non-zeros
  .ROW_PTRS(88'hd0bea6957d6c543f2a1500) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
