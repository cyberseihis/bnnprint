
















module gasId_tnn1_tnnpaar #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 26752'h04180437041404360412042f040a042d040e042a040c0429040604230409042003f1041703f5041503e3040f03ed040d03e5040b03fa040803e4040703da040503d9040403e7040303b9040203cf040103e2040003c403fe03dc03fd03dd03fc03bf03fb03df03f903de03f803ba03f703d503f603bb03f403d403f303c903f203d203f003ce03ef03cc03ee03d103ec03ab03eb03b403ea039303e903c103e803b503e603b003e103a403e003c303db03a003d8038803d703af03d603cb03d3039e03d003bd03cd03a603ca03a903c803a303c703ac03c6038f03c503b103c2038e03c003b703be039503bc03a703b8037c03b6039003b3039403b2038303ae038c03ad033a03aa038103a8038603a5034a03a2036303a10368039f038b039d0364039c0361039b0378039a036903990374039803750397038a039603790392037a0391036f038d0362038903660387035e038503770384036c0382036503800349037f0371037e0306037d034d037b033503760351037303600372033e0370035f036e0359036d0327036b0311036a034403670356035d0333035c0337035b0338035a031c0358032b03570316035502f80354031d03530323035202ff03500345034f033b034e0331034c0307034b0334034802d40347032e034602fa034303360342032f034102dd0340031f033f0328033d0324033c02ef033902fd0332032c03300317032d02f4032a0301032903040326031b03250313032202f7032102d90320030c031e0308031a0315031902ee031802ca031402a8031202c5031002f1030f02e1030e02e6030d02f6030b02f5030a02cf030902d3030502f0030302eb030202b50300025902fe02ce02fc02ec02fb02b002f902e302f3028f02f202c602ed029b02ea02bc02e902cc02e8028802e7028c02e502d002e4028d02e202c702e002da02df02c402de02af02dc02a502db02c202d802b402d7026f02d602b102d502b802d202bd02d102c302cd02bb02cb029e02c902a602c802ab02c1027602c0025702bf02ad02be029a02ba027f02b9029d02b702a902b602aa02b3029202b202a402ae028a02ac029302a7026a02a3029502a2021902a1029902a0026e029f026d029c025a0298028e0297024e02960258029402750291023b02900260028b0279028902020287025c028602300285027d0284027e0283026602820256028101f002800274027c0267027b0247027a0261027802450277025b0273024c027202650271025502700263026c022c026b025d0269025f02680243026402520262022e025e024f0254021c025302460251023e025001f7024d021e024b023a024a02400249020502480219024402370242022702410224023f021f023d0206023c0223023902040238021e023601e4023502310234022f0233022802320200022d0227022b0224022a020802290220022802250226022002260214022502160223021d0222020a022202180221021502210212021f0217021d01d6021c0210021b01e8021b020a02180216021701ed02150213021401fe02130210021201ee021101df021101e9020f01e1020f01ec020c01e5020c0205020901f4020901da020801f6020701d80207019b020601d7020401ff020201ef020101ec020101ff020001f901fe01f901fa01cd01fa01f301f701d901f601f101f4018801f301e001f101de01f001d701ef018701ee01d001ed01e501eb01c101eb01de01e901e301e801da01e7018d01e701dd01e401d201e3019801e101a001e001b001df01d001dd01cc01dc01bd01dc01c001d901b301d8012001d601c601d5019d01d501b801d4016501d401b801d3016c01d301cd01d2014101cc01b001c601bd01c401bc01c4018c01c101ac01c001b201be019101be01bb01bc017501bb01ad01b5016301b5017901b3018901b201a601b1012401b101ad01ae011b01ae019601ac01a701a8019601a8019701a7019c01a601a301a4019d01a4019301a3019601a00165019c0170019b0193019a0185019a01920195012b019401720193015e01900181018f017f018e0169018b0176018a017e01860145018401780183017c0182016e01800140017d0156017b0150017a01130177016c01740136017400ff017401610173016d01710168016f0131016b012e016b015a016a015b01660142016301610162014701600110015e0158015d012f015c0158015a00690156014c0155014e014f0116014f0143014d0116014d012b014c0140014a010e014401050144013801410135014101090141012501400134013c01140139013201370130013701240136012a0135005a013301230132011e0132010a01300128012e0129012d008e012500e801230111012100de011c0117011a00c0011a0107011800da0118010f0116011001150109010f009b010e0100010d0104010900f001080069010800aa01030073010300f6010200fd00fe00a400fd00f100fc008200fb00f300f900f200f800f000f8009a00ee008d00ee00ea00ed00cf00ec00c700ec00d900e800d600e700e100e600d800e500d000e000d700df00b200d9008300d600bc00d500a600d4007b00d400cc00d300b700cd00a000cd007200cb007000ca00bd00c4006800c1009400b800a000b600b300b500ab00b5002100b2009a00b1006400ac00a400a7009500a6009900a3007800a3009c00a2007a00a00051009c0099009b00760099004f0097005300950021009300860091007300900078008d0082008b000f008a001b0085007b00810067007e006a007d0072007c00610079006c007700130074005c0072005a0070002c0070006e006f002d006e00660068001a00600008005f004c005d003e005b000c005900310058000d0057000700560034005500140052000d0050001c004c003a004b0047004900090049003b004600420043002e003f001e0038002f00350022002a00270029000e001f001200190011001800060015000800100005000b01f5021a01ab020e01c7020d01c5020b01970203019f01fd019501fc01c801fb01a501f801a901f201d101ea018a01e601b601e201aa01db01a201cf017c01ce01b701cb011401ca00f401c9018c01c3019e01c201a101bf012001ba016c01b9015401b4008701af0192019901670198018e01940122019100620190008f018f00a1018d0176018b0135018900e9018800230187002c0186017e01850126018400ad018300d1018200fa0181010e01800133017f013c017d0090017b0153017a016f01790040017800360177016401750152017300b90172009e017100fc01700134016b0159016700790165006501640128016300ae01610143015f011b015f0041015e01010157013a0155002b0155008801500074014e0138014b0000014a000701490004014500db014400fb013e010c013900c5012c0032012a010b012900cc0123011d01220014011e003301130063010d00c0010c00c301090101010700b301070084010600e2010400af00ff00e000f800b900ee00d300ed00c200eb00ba00dd007800dc00b800d8000900d7004400d6009400ce007f00ce001300cb00c900ca006b00c8002000c1009700bf00a900bd009600bc00b400bb008300b5009c00b1001000a5003d00a4006f00a1001d009b00380099000e0093008e0092003b008c00480082003d0082007600810068007e0055007d002a007c00300077000300600051005f0045005c00440054004d005300460052003f0051002d004700290039000b0035001c003200210031001f002c001500280019001b0002000f0105016e014e016d0159016a013f0169015401680156016600240162015301600110015d00b0015c0151015a014a0158010f0157000c0152014401510117015000ea01480141014701020147007a0146003c013d00c1013b00e8012d00d4012701000103006100ed00e100e9005e00cf009b00c800b600be004e00ab001300aa005a00a00022009400160085001a00830032006d003a0067003000580017002d001d00250001002000b4015b0119014f0140014d0145014c0074014b01480149013b0146006501430041013f0139013d0012013c00b0013500f200fa000400d2001000bc007200ac00610089002c0069002400310134013e003c013a000201380012013300a001320081012d00d900f8001400da006000680018005a013001420128013700a801360110012e0122012a000901290098012700940123002800f100f901310109012f011e012c0001012b0099012600e9012000d2011b0117011900ca010f00f300fc00db00f400e000e800c500dc003400d8002a00d00084008900920125011601240113011d003b011400bb010e00cc010c0054010700b300d3006a00d1005900c1005b007900930121011a011c000001180052010d00040105005c00f000900091000300410111011f0080011500cb010b0050010300e400ec007000e10043009a001c007c007100730063006b00220062010a01120033010800420106002b010200c200c800c000c40088008c00530074004a004b004000440013001b00c9010400fb0101005100ea001a00c3009c00a30023004900110019007b010000aa00e20048004c000a000b00e300eb000c00a2008a008b000800ab0064006c ;
localparam YMAP = 640'h041d03ff0427042604300434044104380425044004430413041a0431041e041b043a0439041f043b042b043c041c0422043e0435041104190424043204280433043d0442042e04160410043f0421042c;
localparam ADDCNT = $bits(PAAR0) / 32;
localparam FULLCNT = ADDCNT + (FEAT_CNT * 2);
localparam Weights1 = 240'b000100000000000000010000000000000000000010000000000000010100000000010001000100000000000000100000000000000000000000000000000000010011010000000000000000000000000000100000000100000010000100100001000000000000010000100000000010000000010100000000 ;
localparam WNNZ = 240'b000100000000001001110010001000000101100010010000000000010110000000010001001100000000000000100000000000100001000000000000000011010011011000000010000100100100000100100000100100000010100100101111000000011000010110100100010010000100010100000100;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
wire [SUM_BITS-1:0] scorarr [CLASS_CNT-1:0];
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[FEAT_CNT+i] = -feature_array[i];
endgenerate

integer j;
generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam op1 = PAAR0[i*32+:16];
    localparam op2 = PAAR0[i*32+16+:16];
    localparam nodeloc = (2 * FEAT_CNT) + i;
    assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    assign hidden[i] = node[YMAP[i*16+:16]] >= 0;
end
endgenerate

function [7:0] zerocnt(input integer k);
    integer i,j;
    reg [HIDDEN_CNT-1:0] neur1;
    begin
        i = 0;
        neur1 = WNNZ[k*HIDDEN_CNT+:HIDDEN_CNT];
        for(j=0;j<HIDDEN_CNT;j=j+1)
            i = i + !(neur1[j]);
        zerocnt = i;
    end
endfunction

function [7:0] minzc(input integer k);
    integer i,j,h;
    begin
        i = HIDDEN_CNT;
        for(j=0;j<CLASS_CNT;j=j+1) begin
            h = zerocnt(j);
            if(h<i)
                i = h;
        end
        minzc = i;
    end
endfunction

localparam MINZC = minzc(0);

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    localparam Wuse = WNNZ[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wuse[j]) begin
            if(Wneur[j])
                tmpscore = tmpscore + hidden[j];
            else 
                tmpscore = tmpscore + hidden_n[j];
        end
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = 2*tmpscore + zerocnt(i) - MINZC;
    /* assign scorarr[i] = 2*tmpscore + zerocnt(i) - MINZC; */
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
