











module gasId_tnn1_tnnseq #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnn #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(5120'b00000010000000000000000000000000000001000000000000000000000000001000000010000001000000100000000000000000000000001100000000001100000010101000101000000110001010110000010000011010101010110010010100101010000000000010001010000000000000100000000000000110000110101001001000100001000000100000000000000001010000000100000001000000000000000000000000000100000000000110000000000000000000000000100010000000010000000000000000000000000000000000000000000000000011000001101010111010001000110111001100001100000010101010001000110001000010100000100000100000100000100000001000010010000001000000001010100010001100010000101010101000101000011100000001010000010110000000000000000000001000000000000001000100000000000000000000000000000000010000010000000000000000100100000010000000000000000100010100011010101010110011010010101010000101100000101010001000100001100010000100010011001011000000100000000100000000010001000100010100000001010000000000000000000000010000010001000100010000001100010100000000000000000000000010000000110001000000000000000000000001000000000000000000000000000000000011000000011100001000000001000101000110101010101100110100100010110001010000001010100010000000011001100011000100010011110000001100000001100010000100010001000011000001000100000000101000000000001110000100000010000100000001000100000001100000000000000000000000000000000100000000011000000000000001000000000000000000000000000000000000000000000001000000000101100001110010010001000010000110000000000110000110001000001000100000100000101010001010000000000101001000000011000100001000100000001000100010001000010001100010000000000000000000001011000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000100000000000000000000110000000010000001000000110000100111000100001000000011000000001010100010101000010110111010100000000000101100001000101011000101001010011000000010110000110011000101011110100000000000000011000010011100010001110000010000000000000000000000000000000000000000000000000100000000000000100001000000000000000000000000000000100000000000010001001100000000111000101000010110010011010000010000001010101010000000011000100111000001000000101010001000000001100010011100001100001010101000100000000110011001110000110000100011110010100001011000001101000000100000000000000000100000000100000000000000000000000000000100001000000001000000000000000000000100000000000001000000010011100000000111001010010101100000100101001110000000011000100000010110000000010000111000000011100010100001011000000001100111001000110110010000000011100010000101001100000000011001100011010110000000010000000000000000000000000000000001001100000000000000000000000000000000001000000000001100000100000000000010000000000000000001110000001000100110010000000000000000000101000001101010101001000000000010001000000000000000000010000000000000110001000000000000000000000000000000011000000000010000001000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000100000000000000000000010000100000000000000000000000001000000000000100010110000000100000000100100000100000110000001010101000110010010000101010001000100000001011000000100000000000010000001010010000000000001010000100000001001000000000000000000001001100000001000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000001000000000100001001000000101000000001100010000000100000111001000000100000000010100000110100010100100000100001011100001000000001100000110010000110000100001000000000000000000000000000001100100000000010011100001000000010000000100000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000010001000000001001000000000001000000010011000100000001000010101010101000000001100010111100010010001111000001100000001110011000010000100100000000000000001000010000000000000000010000000001000000000001000000110000100000001000000000000000000000010000000000000000000000000000000000000000000100000000100010000000000000000000000100010101001110000010101000101000000110000011000001010101011000100001110010000110000010101100011010010001100001001010010001110000110000000100101010011100100001000111100000001010000000010001000000000001000100000000000000000010000100000000000100000000000010000000000000010000000000000000010001000000000000000000000000000001000100000011000010100000001000000000100000100101000101000110000100011110110001100110100011000000000000000000010010100110001110001000000001001001100111001000010001110000000001001000000000010001100000000101000000010000000000000000000000000011000000000000000010000000000000000000000010010000000000000000001000000010000000000000001110101110000001010001100111000110011100110010001000010111010100010110101000000110001000100001011101010001010010000000010000100000000001100001000101001000000101110010011000000111010100011100111001000100000010000000000000010000000100000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000101100001011001111010010010100000010000111000000101100110000000011000000001000000000000000010001000000100101100000100001000000000011100101000010100000010011000110000000001110010100001001000000001),
  .MASK(5120'b00000010010000000000010010000000000001000000000001000000000000001000000010000001000000100100001000000000000000001100000010011111100011101000111001001110011010111100010110011111111111110111111110101110000000010010011010000100100000101100000000000111110111111101011001100001000000100000011100001101011011000100010001000000000000000000000000000100000000000110000000000000001000000000100010000000010000000000000000000000000000000000000000000000100011011011111011111010011000111111011110011101100011101110011000111001000010100000101100100000100001100000001011010010000001111000011010100110011101010000101010111111101111011100100101011000011110000000000000000000001000000000000001000100000000000010100000000100000100010000010000010001001001100100000010000100100000001101011111111110111110110111111010101010101101111110101111001110111101111011010110110011011011111100101001110101110100111001100101010111110001010101001100010000001011010100011011010100110000111101011100000000010000000000000010000000110001000000000000000000000001000000000000000100000000000010000011000000011100001000000011010101111111101011101101111110100010111011010111001011110011100111011101110111101110011111111010001110011101111011010110011001001011101101000101010011111111000010111110001110101010000100000111000110000001100000000000000100000000000000000100010000011000000000000001000000000000000000000001100000000000000000000001000000000101100111110011010101011010001110110010000111100111011100001001100010100001101010011010101000000111001000010011000101001001100000011000101110101001010001100110000100011010001000101011000100101000100000000000000000000001001100000000000100001000100100000000000110000000000000000000000000000100000000000010000000110000000010000001000100110010101111010100101000000011011110011110110110111001010110111110110101000011101100101010101111101101011011011101101110110010110011011101011111100100000000110011011011011101011001110000010010011000000000000001000000000000000000001001000100000000000010100001000100000001000000000000000000100000000100010011111101100001111001111100011111010011011010010110001010111011101101111100110111000001011000111111001010010001111011011100101101011011111100111001110111111101111011111110110111110111111011111100101101000000100000000001000000100000000100000000000000000000000000000100001000000001000000000001100000000101000010000011101101011111110111010111101011010111110010100111111111001101011010110100111111000100010011111100110111100011110011111110100001100111111100111111110010001011111011111101111101010101011011100111111111001100110000000000100000000000100000000001001100000000000110000000000000000000001100000000001110011100000000000010000000000000000001110101001000110110011100000000010100100101011011101111101101010100000110001000000000011000000010000000000000110001000000000000100000000001001100011000000000010000001000000010100000000000000010010000000000000000000000000000000000010000000000001001100000000100010000000001000000010000100100000000000010100000011000000010000101011110000100100001000100110000100000110111001111101001111110010010101111001000110000001011000000100000000000010100001010010000000001001010100100010001001000010001001000001001001100010001100100000000100100000000000100000000000000000000000100000000000000000010000000010000000000001001000000100001001000000101000010001110010010000100000111001000100101000111011101110111111111110101011111111111100111100001001111110110110111110110111101000000100100000000000000000001100100000000010111100001001000011000100101000001100000000000100000000000000000000001000000000000000100000000001000000000000000000000000010001000000000010000000000010001000000111001100010000001000000010011000100101001011010111111111100010011111011111111011011001111010101101011111111111111010010100100000000001000001000110001000000000001010110000011010001101101011000110000100000001000000000000000000000010000000000000000000000000001000000000001000100000000100010000000000000000000000100010111101111100011101101111111101111010111001001010111111000100101110110001110000011111111011010110111111001001111110001110101111000100101111011111101100111100111110000111010000000010111000000001001000101000100000010000010000110000000000100000000000010010000000100010000000000000000010001000001000000000000000000000001001100101011110110100001111000001010110100100111010101111111000101011110111111101111100011110001000000100110010011111110001111001011000001011011111111101001110001110100001101011011000001110011100110010101010000010001000000000000000000000011000100010000000110000000010000000000000010010000000000000000001000000010010000010000001111111110111011111011100111110110111110110110101011111111110111011111111010111110011100101111111111011101110111001011110010100000101011101001010101101110100111110111011011111111110101011111111011001100000010001000000100010000000100000000000000000000000000100000000000000001000000000000100100000000000100000010000000000100100101101001111011111010011011100011110010111000000101110110100000011100001101000000100011000011001000100110101100000110011000001001011100101010011101010010011011110101010101111010110001101000100001),
  .NONZERO_CNT(640'h3427422822283d33363239252b30332a24333d3328233544252e372f1f3d392639323e2d2d261429),
  .SPARSE_VALS2(58'b1000100000101101101100001111000000101101100010010010010110),  // Bits of not-zeroes
  .COL_INDICES(464'h2419161514110d06040327241816150c0805041d110c2322201d1c1a19110c090600251f1c1513100d0b0a0908002722201f1d1a16130e0a0802), // Column of non-zeros
  .ROW_PTRS(56'h3a302724180c00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
