
















module gasId_bnn1_bnnpaarter #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 59712'h04ef05330001050e05320001051b0531000104d9053000010473052f00010509052e00010510052d00010503052c00010504052b000104db052a000105050529000104ff05280001050205270001050a0526000104ba0525000104ea0524000104f60523000105120522000104fe0521000104c505200001050d051f000104c6051e000104cf051d000104f1051c00010506051a0001046e0519000104f80518000104f90517000104f70516000104e40515000105010514000104fc05130001050f0511000104fb050c00010508050b000104ce0507000104fa0500000104ee04fd000104f204f5000104f304f4000104ac04f0000004ca04ed000004a404ec000004b104eb000004ae04e9000004a604e8000004b504e7000004a204e6000004be04e5000004ad04e3000004ab04e2000004bb04e10000049d04e00000048c04df000004aa04de0000047b04dd0000048404dc0000047504da0000048b04d80000047f04d70000048004d6000004a004d50000049e04d4000004a304d30000048e04d20000048304d10000048f04d00000047604cd0000049304cc0000049c04cb000004af04c90000046d04c80000049504c70000046504c40000047804c30000047004c20000044f04c10000045204c00000046204bf0000046104bd0000043d04bc0000045a04b90000045f04b80000045b04b70000048604b60000041f04b40000043304b30000043f04b20000046004b00000042004a90000042b04a80000042304a70000047904a50000044104a100000485049f00000443049b0000046a049a0000046f04990000048804980000043e04970000041c04960000044804940000042c0492000004070491000003f3049000000428048d000003df048a0000041704890000044a048700000414048200000471048100000446047e00000457047d000003cb047c00000437047a00000451047700000430047400000427047200000449046c000003b6046b0000043504690000041a04680000043c04670000042d0466000004310464000003ff0463000003f9045e0000041b045d00000379045c000003ab04590000041e04580000040a0456000003b00455000003dc045400000432045300000419045000000415044e0000040e044d000003d0044c000003f4044b000004050447000003be0445000003ce0444000004110442000004100440000003d7043b0000042a043a000003e80439000004020438000003c2043600000354043400000412042f000003f0042e000003ca0429000003ec0426000003970425000003e604240000038d04220000039c0421000003ed041d000003fa0418000003480416000003b5041300000367040f000003ac040d000003c5040c000003da040b0000035b04090000033004080000038f0406000003cd0404000003b10403000003860401000003de0400000003cc03fe000003db03fd000003bb03fc000003ae03fb0000039903f8000003bc03f7000003c103f6000003e303f5000003d503f2000003d203f10000038e03ef000003c703ee000003bd03eb000003c803ea000003d603e90000038903e7000003a703e50000034e03e40000037703e2000003a303e1000003b803e0000003c003dd0000036203d90000036d03d80000034303d4000003a103d30000037e03d10000037103cf0000030103c90000037203c60000037f03c40000036003c30000036a03bf0000038303ba0000039a03b9000002b503b70000032b03b40000031703b30000039403b20000039e03af0000033603ad0000037b03aa0000036c03a90000030a03a80000039203a60000037a03a50000036803a40000037603a20000038403a0000002de039f0000037c039d0000033a039b000002f103980000032503960000038003950000035903930000035f0391000003700390000002dd038c00000334038b0000034a038a000003190388000003200387000002f603850000035e038200000361038100000347037d000002ea03780000036f03750000030003740000034903730000031a036e00000329036b0000033803690000031f03660000034f0365000002ef0364000002d00363000002e3035d00000323035c000002e5035a000002e803580000032d0357000002fb0356000003120355000003260353000002e40352000002d40351000002af035000000316034d0000030d034c0000030e034b0000030c0346000003070345000003020344000002fa0342000002ce034100000278034000000327033f000002d2033e00000306033d000002e7033c00000313033b000002fe0339000003090337000002ed0335000002bd0333000002e60332000003220331000002fc032f0000031e032e0000030f032c000002ee032a000003150328000002eb0324000003080321000002c4031d000002c2031c000002a6031b000002520318000002ba0314000002620311000002e00310000002f7030b000002d50305000002f20304000002ec0303000002c702ff0000027f02fd0000028402f9000002c802f8000002bc02f50000027e02f40000025502f3000002ac02f0000002d302e90000026c02e20000028102e1000002c502df000002a302dc0000023a02db000002aa02da000002c902d9000001dc02d8000002cd02d7000002b802d60000027102d10000029e02cf0000027902cc000002b402cb000002ab02ca0000023202c60000029502c30000027002c10000028a02c00000028302bf0000026602be0000027a02bb0000020902b90000027702b70000026002b60000027d02b30000027102b20000027602b10000022b02b0000001cc02ae0000029902ad0000022802a9000001c002a80000029302a70000025902a50000028602a40000024602a20000027c02a10000029b02a000000289029f0000027b029d0000028f029c0000027a029a0000022e02980000028802970000022402960000027902940000028d029200000274029100000270029000000275028e00000273028c0000027c028b0000024602870000026e0285000002580282000001ea02820000022d028100000256028000000254027f0000026f027e00000263027d00000247027800000225027700000236027500000256027300000258027200000221027200000239026f00000269026e0000025e026d00000227026c00000268026b0000023e026b0000025a026a000002180269000001cd02680000023402670000022f02670000023c02660000026102650000026102640000025d02640000022d025f000001f8025e00000242025d0000024d025c00000221025c00000225025a000001fc02590000025002570000024202570000015f0255000001f902530000021e02520000024402510000023a02510000020a02500000020b024e000001ba024e00000107024d0000024a024b000001e2024b0000018b024a000001aa02490000017e02490000021d02480000021202480000023302470000021b0244000000f502410000022f0240000001fe02400000021f023f0000021e023f00000223023e000001da023c0000022b02390000022c0238000002190238000001fd0236000001ba02340000020e0233000002170232000002280231000001a8022c000001e2022a0000021a0229000002020229000001fe02270000020e0226000002000224000001ab02220000020c0220000001de021d00000196021b000001f5021a000002100218000001b102170000020602160000019c0216000001d40213000001b50213000001720212000002050211000001b70210000001db020c00000205020b000001c8020a000002060209000001db0208000001cc0208000002010202000001590201000001cd0200000001ad01fd000001d901fc000001ae01fb0000018001fb0000019e01fa0000017c01fa000001cb01f9000001e101f8000001e601f7000001d501f7000001ec01f6000001eb01f6000001d801f5000001a301f4000001cd01f0000001c701f0000001e701ef000001c201ee0000018d01ee000001b301ed000001d401ec000001e601eb0000018201ea000001e501e8000000e301e7000001e401e50000014d01e4000001cf01e1000001d801e00000010c01e0000001d201df0000017e01de0000012001da000001d201d7000001c101d7000001d101d6000001bb01d6000001b201ce000001ad01ce000001bf01cb0000019d01cb0000019a01ca0000019a01c9000001be01c7000001ae01c60000014401c5000001ba01c40000017401c3000001b001c1000001ad01bd0000017601bc0000019a01b90000019d01b80000019001b70000016001b70000017e01b60000018301b50000011f01b40000016701af0000018701ac0000019001a80000016501a80000016201a70000018501a60000019401a50000019901a20000016e01a000000139019f00000177019d0000014a019b0000018e01980000017301970000014e0197000000f901970000019201960000018101960000018901950000014201940000016f019300000155019100000183019000000137018d00000154018b0000015c01890000015b01880000014801880000013901860000017101850000013f01840000017001820000015e018100000156018000000177017f0000011f017f00000155017c00000146017a00000120017500000169017100000161017000000156016f000000fc016b00000167016a0000014a0169000000b10168000000890168000001420166000001370165000001470164000000ee0161000000e60160000000e9015d0000015a015c00000133015c0000014501580000010c0158000001530157000000c401550000013e0154000001410152000001490151000000d9014f0000012a014d00000104014c000000ab014c00000126014b000001470148000001320146000001300146000000de01430000013c014100000124013e00000120013e00000110013d00000110013b0000012801360000011d01360000011b01360000011601360000011a01350000011401350000012e0131000000ab013100000118012f00000121012b000000ff012b000001240127000000e00123000000c901230000010201220000010c011f000000dc011e00000115011b000000bd011a000001010119000000d601180000010d0117000001070114000001000114000000e80113000000890112000000810111000000fc010e000000f9010e00000102010c000001060107000000f60106000000ec0106000000f401050000009c0102000000fb0101000000cc0101000000ef0100000000ce00ff000000a900ff000000e500fe000000d000fc000000f800fb000000f400f80000009a00f7000000ed00f6000000dc00f40000009100f2000000ec00f1000000bf00f00000009200ef000000dd00ee0000009c00e8000000dd00e6000000de00e4000000b500e20000009000e1000000d400df000000c800dc000000d700da000000be00da000000b400da000000cd00d9000000d500d8000000cf00d5000000a600d30000009500d20000009100d20000008f00d10000008d00d10000008d00d00000009700ce000000a900cc000000b100cb0000008d00cb000000b400c7000000bf00c2000000a300c0000000b900bb000000ac00ba000000a100b9000000a700b80000009600b80000008400b70000002400b7000000aa00b3000000ac00b20000008700b20000008f00ae000000a500ab0000009800aa0000008800a70000009800a60000009b009f0000009400990000007c00800000026a027b000100ec02760001012a0262000102530254000100df022e0001016402190001019401d5000100ee01c7000100d20173000100bd0128000100f102800000010502740000014e026d000001e80265000001230263000000b50260000000de025f000001cc0241000000f80231000000aa022a0000011702260000021f0223000001c10222000001dc0220000001d102110000011f01f4000001ce01ef0000015d01ed0000017401df0000014901d90000017e01b50000014d01ae000000d10190000000fb0131000001af025b00010122024f000100b3024c000101bf02450001019202430001002b023d000101890237000101bb0215000100d60204000100ea01ff000101b301f20001016c01f10001010901d30001013501cf0001008401ca000101a701b9000100d001b1000100db019b0001017f019900010163019800010153019500010094018a000100b80157000101180150000100900142000100af01380001010e012e000100a9012d0001009b012c000100cf0128000100eb0125000100f20124000100ef012100010016011c000100c400f200010064006c000101f3023b000001d002350000018f0230000001bc021c0000017d02140000019f020f000001b6020d000001ac0207000001790203000000b101e9000001c901e30000014f01dd0000018301c8000000cd01c60000012601c5000001a501c4000000ab01c3000001a001c20000013701c0000001ab01be000000e801bd0000013f01b8000000ad01b40000015e01b2000000cd01b00000014b01aa000000ba01a3000000c701a200000141019e000000d7019c000001410193000001670191000000f4018f00000023018d0000016d018c00000119018b00000080018a0000015c01880000015f018500000110018100000125018000000089017d00000159017b000000c0017b0000013d0179000000c80177000001440174000000f1017300000100016f000000e1016d000000d101650000014201640000011e0163000000eb01610000010b015b000000e0015b0000011f015a000000e901590000008b0155000000d30152000000f80151000000d6015100000112014f0000013a014b000000ac0146000001270145000000a40145000000900144000000b30143000000e40140000000c101400000009e01400000009501390000012701360000010f0134000000bb0133000000f70132000000e70130000000e7012d000000af012b000000e2012a000000d40129000000bb0129000000ed011d000000bc011b000000ce0119000000cc0116000000880115000000a601140000008701130000009a0110000000f90108000000c60108000000aa0107000000810104000000d80103000000c70100000000be00fe000000d400fd0000009e00fa000000e100f50000009d00f0000000b900e5000000c900e20000009a00e00000009f00dc000000cf00d9000000be00d9000000c300ce0000000300c90000002400c6000000a700c20000009d00b9000000880092000001270182000101130171000100fb0169000100e80153000100dd015200010094014d000100ad013500010112011d000100b500e2000100ad00da0001009200cb000100a600c0000100eb01a6000000ae018c0000015a017c0000011f01700000015e01680000013c015f000000890157000000ff0143000000b70137000000a5012d000000cb010e000000f80105000000e301050000008b00f2000000de00e200000095013900010003016c0000009b00ec0001008601a90001007b01a100010184018e0001014e017a000100dc01750001012b016e0001009401660001015401600001014a015d000100c40158000101170148000100d8013c000100d70133000100ff012e000100e3010f0001009900e70001008c00c6000100a000b00001010201a40000016a0187000001560186000000fe017600000147016b000000a90150000000b70149000000b2013f0000010a013e00000096013d000000b4012a000000e80128000000c5011a000000d80119000000f10117000000bf0115000000fc011000000097010a000000870101000000b100fa000000bc00f70000009700e1000000d300e00000009200db000000a200c7000000c000c30000002e0093000000530073000000ff0172000101300162000100f9011d000100c1011a000100a40104000100d200e90001010e014c000000d00132000000980131000000f401290000012401250000010d0111000000c500ef000000ab00e3000000aa00d30000008901150001009f0126000000f0010b0001010b01180000007c008f000000a5017800010084013a00010109012c000101120122000100e5011b000100b60109000100b00103000100b400f8000100b300f60001009000f50001009d00ee000100a000ea000100dd00e2000100d900db0001009c00ba000100530082000100a80138000000bd0134000000240123000000c40121000000b20114000000be010f000000d1010a000000bf0104000000e401010000009900fd000000e600ed000000da00e3000000ae00cb000000b800ca0000008800b70000008600a8000000120043000000c50113000100a20102000100a300f9000100d200f4000100b100b5000100960120000000a10105000000c100e8000000d500d70000008b0095000100b001030000009100f7000100ce00de000100de00fe0000009e0100000000c9012f000100cd011e000100b5010c0001008900cf0001009c00cc0001000300830001002e011100000093010d0000009a0107000000fc00fd0000008c00f5000000ef00f3000000df00f2000000b900f10000008d00ed000000d500d6000000bc00d40000001a004b000000c700f60001009e00c60001008f013b000000a900c3000000a600ba0000009700f0000100ae00e10001009d00ee0000008600fa000000bc0108000100b200fb000100e70116000100d500e4000100af00e00001009f00a20001007c008500010049006300010000004200010008000c00010016011c000000a000ea000000e500e90000009800ca0000009100ac00000024008a000000100041000000b300eb000100be00db0001009900b40001009400d9000000c000ec000100df00e6000100ad00bb00010051007900010040004400010022002a000100d80106000000d400dc000000d200d6000000a300a7000000dd00f3000000d700da000100b800c1000100ce00d300010034006b00010019001b0001000a000b000100c800cf0000009b00b600000027005500000006004f000000ab00d1000100a500c1000100a100a40001003b00740001001c006a0001001100590001001e005800010048004a0001002100620000000200280000002e00cd0000009200c700000016008e00010052007000010013003d0001005c00750000002d006e00000036006600000017006500000001005a0000003f0056000000050045000000200029000000c600cc000000bc00d0000100600068000100c900ca0000003a007d0000003700770000000900690000001800570000002c004c0000000d0025000000c800cb0001005f007f0001005b00710001005d006f00010031004d0001002f003c000100be00c000000015007800000061007200000032006d0000001d006700000038005e0000000700350000001f0033000000ab00c5000000300050000100460047000100b800c40000003900540000000e0014000000b300b4000100a500b20000000f007e0001000400760001009200b50000003e004e000000ad00bb000000ba00c3000100a100a40000009e00ae0000009b00b6000100a000b00000009d00b90001009f00a2000000a900b100010026007a0000009400bf0001009900b7000100a300a7000100a600af0000009100ac00010097009c0001008900980000008600a80001008f00aa0000009a00bd0000009500c200000016008e00000026007a0001002e00930001009000960000008c008d00010088008b0000003e004e0001000f007e0000000400760000000e001400010024008a0001003000500000004600470000003900540001006100720001005b00710000001500780001001d006700010038005e0001005f007f0000005d006f00000031004d0000002f003c0000000700350001008400870000001f003300010032006d0001000d00250001006000680000007c00850000003a007d0001000900690001001800570001002c004c0001003700770001001700650001005c007500010036006600010001005a0001003f00560001000500450001002000290001002d006e00010052007000000013003d0000003b00740000002100620001000300830000001c006a00000011005900000048004a0000000200280001001e005800000027005500010006004f00010019001b00000034006b0000000a000b00000022002a00000051007900000040004400000053008200000010004100010000004200000049006300000008000c0000008000810000001a004b00010012004300010073007b00000023002b00000064006c0000 ;
localparam YMAP = 1280'h000005360000053e00010538000005540000055a00010545000005460000055200010558000005420000053b000005500001053d000105430000055500000557000005390001055900000549000105340001054e000105400001054f00000537000005510000053a000005530000055b0001053f000105470001055600000541000105350001054a0000053c0000054b0001054c0000054d0000054400010548;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 240'b001101100010110011101111111110000101100100111011101110001100100011010110111110010011010000101000111011101111100011011101110101110110000001111111010010111010101110110110000010000111110101011111100011100111010010101100110110001100101001011011 ;
localparam WIDTH = 320'h09090909090909090a0909090a080a09090809090908080909090a0808090909080808080a080909;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;
generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam subad = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(subad)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] < 0;
    initial begin
        #20
        $display("%b, %d | %d", signy, ymap, node[ymap]);
    end
end
endgenerate

initial begin
    #10
    for(j=0;j<FULLCNT;j=j+1) begin
        $display("%d | %d | %b, %d, %d", j, node[j], PAAR0[(j- FEAT_CNT )*48],  PAAR0[(j-FEAT_CNT)*48+16+:16], PAAR0[(j-FEAT_CNT)*48+32+:16]);
    end
end

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wneur[j])
            tmpscore = tmpscore + hidden[j];
        else 
            tmpscore = tmpscore + hidden_n[j];
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = tmpscore;
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
