module xnorpop (input [15:0]a, output [49:0]o);
assign o[4:0] = !a[0] + a[1] + !a[2] + a[3] + a[4] + a[5] + !a[6] + !a[7] + !a[8] + !a[9] + !a[10] + !a[11] + !a[12] + a[13] + !a[14] + !a[15];
assign o[9:5] = a[0] + !a[1] + !a[2] + a[3] + a[4] + !a[5] + !a[6] + !a[7] + !a[8] + a[9] + a[10] + a[11] + a[12] + !a[13] + a[14] + !a[15];
assign o[14:10] = !a[0] + !a[1] + !a[2] + !a[3] + !a[4] + !a[5] + !a[6] + a[7] + a[8] + !a[9] + a[10] + a[11] + !a[12] + !a[13] + a[14] + !a[15];
assign o[19:15] = !a[0] + !a[1] + a[2] + a[3] + !a[4] + !a[5] + a[6] + !a[7] + !a[8] + !a[9] + !a[10] + a[11] + !a[12] + !a[13] + !a[14] + a[15];
assign o[24:20] = !a[0] + a[1] + a[2] + !a[3] + !a[4] + !a[5] + a[6] + !a[7] + a[8] + !a[9] + a[10] + !a[11] + a[12] + a[13] + a[14] + !a[15];
assign o[29:25] = !a[0] + !a[1] + a[2] + !a[3] + a[4] + a[5] + a[6] + a[7] + a[8] + a[9] + a[10] + !a[11] + !a[12] + a[13] + !a[14] + a[15];
assign o[34:30] = a[0] + a[1] + !a[2] + !a[3] + a[4] + !a[5] + a[6] + a[7] + a[8] + a[9] + !a[10] + a[11] + !a[12] + !a[13] + !a[14] + !a[15];
assign o[39:35] = !a[0] + !a[1] + a[2] + !a[3] + !a[4] + a[5] + !a[6] + a[7] + !a[8] + a[9] + a[10] + a[11] + a[12] + !a[13] + !a[14] + !a[15];
assign o[44:40] = !a[0] + !a[1] + a[2] + a[3] + a[4] + !a[5] + !a[6] + a[7] + !a[8] + a[9] + !a[10] + !a[11] + !a[12] + a[13] + a[14] + !a[15];
assign o[49:45] = !a[0] + a[1] + !a[2] + a[3] + a[4] + !a[5] + a[6] + !a[7] + !a[8] + a[9] + a[10] + !a[11] + !a[12] + !a[13] + a[14] + a[15];
endmodule
