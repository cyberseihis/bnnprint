module seqq #(
  parameter N = 4,
  parameter B = 4,
  parameter M = 4
  ) (
  input clk,
  input rst,
  input [N*B-1:0] data,
  output [M-1:0] out
  );
  
  reg [$clog2(N)-1:0] cnt;
  wire [M*N-1:0] weis;
  wire [M-1:0] weit;
  wire [B-1:0] in;
  wire put;
  
  assign weis =
      `include "weis.wei"
      ;
  genvar i;
  generate
    for (i=0;i<M;i=i+1) begin
      accum #(.N(N), .B(B)) acc1 (
        .data_in(in),
        .clk(clk),
        .put(put),
        .rst(rst),
        .add_sub(weit[i]),
        .out(out[i])
      );
    end
  endgenerate

  assign put = cnt==N-1;
  assign in = data[cnt*B+:B];
  assign weit = weis[cnt*M+:M];

  always @(posedge clk or posedge rst) begin
      if(rst || cnt == N-1) begin
          cnt <= 0;
      end
      else begin
          cnt <= cnt + 1;
      end
  end
  
endmodule
