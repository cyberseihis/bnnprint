
















module winered_tnn1_tnnpaarter #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 5424'h0009005d00010016005c0001000a005a0001003f005800010004005700010001005300010011005000010034004f00010000004e00010001004d00010006004c0001000900490001000d00480001003b00470001001900440001002500430001003900420001000700410001001d00400001002c003c0001003200370001002b00330001001c002f0001001c002e0001000b00280001000900260001002300240001000f002300010029004b0000001c004600000020004500000021003d0000001a003a0000002200380000001600360000003000350000000d003100000018002d00000004002b0000000b002a00000009002a0000001200290000001a00280000001000270000000300270000002400260000001900250000001e002100000006002000000011001f0000000b001f0000001d001e00000005001b00000004001b00000014001a0000000b00180000001500160000000600150000000100150000000800140000001000130000000900120000000700100000000d000f00000000000f0000000d000e00000002000e00000001000c0000000700090000000500090000000600080000000100050000000000030000000000020000000c00220001000000030001000f001b0000000100190000000e00150000000600100000001100180001000a001700010004001700010002001300010007000e00010008000b0001000f00140000000c00130000000e001200000003000f00000008000d00000008000a00000002000e00010000000200010004001200000000001000010009001100010001000600010003000a00000005000800010007000c00000001000400000003000d00010000000c00000007000900010003000b00000006000a00010002000500010007000800010000000400000009000a0000000200050000000100060000 ;
localparam YMAP = 1280'h0000006800010060000000160001007400000078000000710001006b000100720000006a0001006500010070000000510001004a0000006c0000006d00000077000100690001005b00000056000100670001006e0001005f0000005e0000007900010062000100520001007b000000760000005400010063000100640001006f000000750000003e000100730000007a00010055000000590000006600010061;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 240'b001010100100001000000000001000000100000000110011000000000100000001001000100001000000001100000000100000000000000001000000000000100000000000000000011000010001000000001000001000000000000000101110000000001000000001010000010000000000000000010100 ;
localparam WNNZ = 240'b001010100100001000000000011100010101000100110011101000100101000011011000100011111000011100000000100000000001000001000010000010100000001000000000011100110001001100001000001100000000000000101110001000001000000001110100110001100001000000011101;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
wire [SUM_BITS-1:0] scorarr [CLASS_CNT-1:0];
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;

generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam adsub = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(adsub)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] <= 0;
end
endgenerate

function [7:0] zerocnt(input integer k);
    integer i,j;
    reg [HIDDEN_CNT-1:0] neur1;
    begin
        i = 0;
        neur1 = WNNZ[k*HIDDEN_CNT+:HIDDEN_CNT];
        for(j=0;j<HIDDEN_CNT;j=j+1)
            i = i + !(neur1[j]);
        zerocnt = i;
    end
endfunction

function [7:0] minzc(input integer k);
    integer i,j,h;
    begin
        i = HIDDEN_CNT;
        for(j=0;j<CLASS_CNT;j=j+1) begin
            h = zerocnt(j);
            if(h<i)
                i = h;
        end
        minzc = i;
    end
endfunction

localparam MINZC = minzc(0);

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    localparam Wuse = WNNZ[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wuse[j]) begin
            if(Wneur[j])
                tmpscore = tmpscore + hidden[j];
            else 
                tmpscore = tmpscore + hidden_n[j];
        end
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = 2*tmpscore + zerocnt(i) - MINZC;
    /* assign scorarr[i] = 2*tmpscore + zerocnt(i) - MINZC; */
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
