
















module winewhite_tnn1_tnnpaarter #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 4848'h000f005200010009005100010038004e00010022004c00010023004b00010011004a00010003004900010009004700010033004500010013004200010011004100010011003e0001002e003c00010037003b0001000f003a0001003200360001001f00350001002000300001002d002f0001000600290001001300270001000200250001000700220001001600210001000600210001000f002000010019001f00010013001c0001001400160001002300400000002b00390000001200340000001c003100000019002c0000000e002a0000000c00280000000700260000000900250000001100240000000100240000000f001e0000000b001e00000010001d00000005001d00000019001c0000000e001b00000005001a0000000800180000000300180000000400170000001500160000001100140000000d00140000000d001300000007001200000000000d0000000000110000000b00100000000300100000000b000e0000000a000e00000006000d00000008000c00000008000b00000001000b00000008000a00000003000a0000000700080000000200060000000f00180000000800140000000a001000000007000d0000000a000c00010008001b0001000b001a0001000500090001000600170000001200150000000000120000000a000f00000003000c0000000100070000000d000f00000004000d0001000900100000000c000e00000002000a00000003000500000002000600010004000e00000003000700000000000100000001000500010006000c00000000000800000006000b00000003000900000005000a0000000100020000000400070000 ;
localparam YMAP = 1280'h0000006000010026000000570000006e000100690001006400010044000100460001005b000100500000006d0000000a0001003d0000003f0000005d000000620001004f0001006c000100670001006100000058000100630000005e000100430000005c000000550000005a0001006b0000006a000100590000005f0000006500000054000100680001005300010066000100560001006f0001004d00000048;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 280'b0010000000000001000101000010000000110000000000001000000000000000000000000000000000000000000100000100000000000000000000000010000010000001100000011000000000000010001100000000000100010100000000000000000001100000000100010101100000001000100000000000000000010000000101001000100010010000 ;
localparam WNNZ = 280'b0110111101001001100101110011000001110110000000101000000010000001001010000000000000000010000100000110000100010001000000000010001010000001100000011000000000000010001100100000001100010100000000100000000001100100110100011101100100001100100000000100000000010000100101011000111011010010;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
wire [SUM_BITS-1:0] scorarr [CLASS_CNT-1:0];
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;

generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam adsub = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(adsub)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] <= 0;
end
endgenerate

function [7:0] zerocnt(input integer k);
    integer i,j;
    reg [HIDDEN_CNT-1:0] neur1;
    begin
        i = 0;
        neur1 = WNNZ[k*HIDDEN_CNT+:HIDDEN_CNT];
        for(j=0;j<HIDDEN_CNT;j=j+1)
            i = i + !(neur1[j]);
        zerocnt = i;
    end
endfunction

function [7:0] minzc(input integer k);
    integer i,j,h;
    begin
        i = HIDDEN_CNT;
        for(j=0;j<CLASS_CNT;j=j+1) begin
            h = zerocnt(j);
            if(h<i)
                i = h;
        end
        minzc = i;
    end
endfunction

localparam MINZC = minzc(0);

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    localparam Wuse = WNNZ[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wuse[j]) begin
            if(Wneur[j])
                tmpscore = tmpscore + hidden[j];
            else 
                tmpscore = tmpscore + hidden_n[j];
        end
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = 2*tmpscore + zerocnt(i) - MINZC;
    /* assign scorarr[i] = 2*tmpscore + zerocnt(i) - MINZC; */
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
