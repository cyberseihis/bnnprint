













module winered_bnn1_bnnroperm #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 440'b00111000000010010101000001100100000010101100111011111111100110010010101011011111011001111000000011011011110000101110011001010100111001100010011111111000001011011000111010100001111000000011111111011001010011110111100100101111100010100101010011011100011010000111000110100000101000001111001010010111010000111110001000001110110011100011111010111001101100001110001100111011110110001110100110001011101101101011101001101010001110111011100110011000 ;
  localparam Weights1 = 240'b101111011011111011101101100111001000110011101100101011111101111011110100000010100110100100101101111011000011011010101101100011010011101001001000010000100010010101111011110010101001100010001101000100010100111010011100001000001001100000110101 ;

  romesh_seq #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
