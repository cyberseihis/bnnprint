`timescale 1us/1ns









module tbHar_bnn1_bnnpar #(

parameter FEAT_CNT = 12,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)();
reg clk;
reg [FEAT_CNT*FEAT_BITS-1:0] features;
wire [$clog2(CLASS_CNT)-1:0] prediction;
wire [FEAT_CNT*FEAT_BITS-1:0] testcases [TEST_CNT-1:0];
parameter Nsperiod=5000;
parameter period = Nsperiod/500;


assign testcases[0] = 48'hb9811498a121;
assign testcases[1] = 48'hb9700187a110;
assign testcases[2] = 48'hb9700088a000;
assign testcases[3] = 48'hb9700088a000;
assign testcases[4] = 48'hb97000889000;
assign testcases[5] = 48'hb97000889000;
assign testcases[6] = 48'hb97000899000;
assign testcases[7] = 48'hb97000889000;
assign testcases[8] = 48'hb97000889000;
assign testcases[9] = 48'hb97000889000;
assign testcases[10] = 48'hb97000889000;
assign testcases[11] = 48'hb97000889000;
assign testcases[12] = 48'hb97000889000;
assign testcases[13] = 48'hb97000889000;
assign testcases[14] = 48'hb97000899000;
assign testcases[15] = 48'hb97000799211;
assign testcases[16] = 48'hb97112888000;
assign testcases[17] = 48'hb97011889000;
assign testcases[18] = 48'hb97000889000;
assign testcases[19] = 48'hb9701088a101;
assign testcases[20] = 48'hb8701188a101;
assign testcases[21] = 48'hb97011899111;
assign testcases[22] = 48'hba8111899123;
assign testcases[23] = 48'hba8011889013;
assign testcases[24] = 48'hb97000889000;
assign testcases[25] = 48'hb97000889000;
assign testcases[26] = 48'hb97000889000;
assign testcases[27] = 48'hb97000889000;
assign testcases[28] = 48'hb97000889000;
assign testcases[29] = 48'hb97000889000;
assign testcases[30] = 48'hb97000889000;
assign testcases[31] = 48'hb9701188a001;
assign testcases[32] = 48'hb9700089a000;
assign testcases[33] = 48'hb97000889000;
assign testcases[34] = 48'hb97000889000;
assign testcases[35] = 48'hb97000889000;
assign testcases[36] = 48'hb97000889000;
assign testcases[37] = 48'hb97000889000;
assign testcases[38] = 48'hb97000889000;
assign testcases[39] = 48'hb97000889000;
assign testcases[40] = 48'hb97000889000;
assign testcases[41] = 48'hb97000889000;
assign testcases[42] = 48'hb97000889000;
assign testcases[43] = 48'hb97000889000;
assign testcases[44] = 48'hba61126a5112;
assign testcases[45] = 48'hb97011797102;
assign testcases[46] = 48'hb97000799001;
assign testcases[47] = 48'hb97000889000;
assign testcases[48] = 48'hb97000889000;
assign testcases[49] = 48'hb9700088a001;
assign testcases[50] = 48'hb9701088a000;
assign testcases[51] = 48'hb87000889000;
assign testcases[52] = 48'hb97000889000;
assign testcases[53] = 48'hb97000899000;
assign testcases[54] = 48'hb97000889000;
assign testcases[55] = 48'ha9710086b111;
assign testcases[56] = 48'hb9700087a011;
assign testcases[57] = 48'hb97000889000;
assign testcases[58] = 48'hb97000889000;
assign testcases[59] = 48'hb97000899000;
assign testcases[60] = 48'hb97000899000;
assign testcases[61] = 48'hb97000899000;
assign testcases[62] = 48'hb97000889000;
assign testcases[63] = 48'hb97000889000;
assign testcases[64] = 48'hb97000889000;
assign testcases[65] = 48'hb97000889000;
assign testcases[66] = 48'hc9721196e102;
assign testcases[67] = 48'hc9710086b112;
assign testcases[68] = 48'hb9700087a001;
assign testcases[69] = 48'hb97000889001;
assign testcases[70] = 48'hb97000889000;
assign testcases[71] = 48'hb97000889000;
assign testcases[72] = 48'hb97000899000;
assign testcases[73] = 48'hb97000889000;
assign testcases[74] = 48'hb97000889000;
assign testcases[75] = 48'hb97000899000;
assign testcases[76] = 48'hb97000889000;
assign testcases[77] = 48'hc97000889000;
assign testcases[78] = 48'hb97000899000;
assign testcases[79] = 48'ha976766b9456;
assign testcases[80] = 48'hb9877679a456;
assign testcases[81] = 48'hc97687889455;
assign testcases[82] = 48'hb97587889455;
assign testcases[83] = 48'hb97577889455;
assign testcases[84] = 48'ha97666889455;
assign testcases[85] = 48'hba7666889456;
assign testcases[86] = 48'hc97676889446;
assign testcases[87] = 48'hc97677899456;
assign testcases[88] = 48'hc97576799555;
assign testcases[89] = 48'ha9767689a556;
assign testcases[90] = 48'ha98677899557;
assign testcases[91] = 48'hc97677899556;
assign testcases[92] = 48'hb97676889555;
assign testcases[93] = 48'haa766687a456;
assign testcases[94] = 48'hb976665c9455;
assign testcases[95] = 48'hc877776a9455;
assign testcases[96] = 48'ha97776799556;
assign testcases[97] = 48'hba867688a555;
assign testcases[98] = 48'hc97676889455;
assign testcases[99] = 48'hb87676889455;
assign testcases[100] = 48'hba7676889555;
assign testcases[101] = 48'hba7676889455;
assign testcases[102] = 48'hc97676889556;
assign testcases[103] = 48'hb87776899556;
assign testcases[104] = 48'ha9767679a455;
assign testcases[105] = 48'hba8677889455;
assign testcases[106] = 48'hc87687899456;
assign testcases[107] = 48'hb87686899455;
assign testcases[108] = 48'hb97577889455;
assign testcases[109] = 48'hc87988799446;
assign testcases[110] = 48'hc96a87799356;
assign testcases[111] = 48'hba89996b9747;
assign testcases[112] = 48'h9989995b9647;
assign testcases[113] = 48'h89799787a557;
assign testcases[114] = 48'hc97aa87a9867;
assign testcases[115] = 48'hba7ba9799877;
assign testcases[116] = 48'hb87baab59568;
assign testcases[117] = 48'hd87a99b69468;
assign testcases[118] = 48'hb96a9a69b466;
assign testcases[119] = 48'hc96b8b79a467;
assign testcases[120] = 48'hd96bad4db878;
assign testcases[121] = 48'ha96bbc69aa78;
assign testcases[122] = 48'haa7bab78aa68;
assign testcases[123] = 48'hb97aac79a978;
assign testcases[124] = 48'hb87cacb77667;
assign testcases[125] = 48'hb98daca67668;
assign testcases[126] = 48'hb87eae4bf758;
assign testcases[127] = 48'hba7b8d3cf868;
assign testcases[128] = 48'hb97a8d5bd97a;
assign testcases[129] = 48'hba8bad89a779;
assign testcases[130] = 48'hd96cbe79a979;
assign testcases[131] = 48'ha87c9e967a69;
assign testcases[132] = 48'ha97badc55667;
assign testcases[133] = 48'hb9379b4b9469;
assign testcases[134] = 48'ha847986b947a;
assign testcases[135] = 48'ha9778898856a;
assign testcases[136] = 48'hba7688b56759;
assign testcases[137] = 48'hb9679a979769;
assign testcases[138] = 48'ha9678889867c;
assign testcases[139] = 48'ha9778798876c;
assign testcases[140] = 48'hba588b6ac66a;
assign testcases[141] = 48'hba578b5bb37a;
assign testcases[142] = 48'h89379c49b56a;
assign testcases[143] = 48'hab378d7aa76b;
assign testcases[144] = 48'hb9678ba9776d;
assign testcases[145] = 48'hb9779ab7575c;
assign testcases[146] = 48'ha977ab99a85b;
assign testcases[147] = 48'hba68ab98876e;
assign testcases[148] = 48'hba779c88987f;
assign testcases[149] = 48'h99778c5bf76b;
assign testcases[150] = 48'h86579c5be65b;
assign testcases[151] = 48'hb9678d7aa74a;
assign testcases[152] = 48'hb9769ba7475f;
assign testcases[153] = 48'hb9769ca7575f;
assign testcases[154] = 48'hb9668c89a74b;
assign testcases[155] = 48'ha9769d98886d;
assign testcases[156] = 48'hb9879e79c87d;
assign testcases[157] = 48'hb8779e5af76a;
assign testcases[158] = 48'ha88114989111;
assign testcases[159] = 48'hb9601088a100;
assign testcases[160] = 48'hb9600088a000;
assign testcases[161] = 48'hb9700188a000;
assign testcases[162] = 48'hb97000899000;
assign testcases[163] = 48'hb97000899000;
assign testcases[164] = 48'hb97000889000;
assign testcases[165] = 48'hb97000889000;
assign testcases[166] = 48'hb97000889000;
assign testcases[167] = 48'hb97000889000;
assign testcases[168] = 48'hb97000889000;
assign testcases[169] = 48'hca8013898001;
assign testcases[170] = 48'hb96000889000;
assign testcases[171] = 48'hb97000889000;
assign testcases[172] = 48'hb97000889000;
assign testcases[173] = 48'hb97000889000;
assign testcases[174] = 48'hb97000889000;
assign testcases[175] = 48'hb97000889000;
assign testcases[176] = 48'hb97000889000;
assign testcases[177] = 48'hb97000889000;
assign testcases[178] = 48'hb97000889000;
assign testcases[179] = 48'hb97000889000;
assign testcases[180] = 48'hb97000899001;
assign testcases[181] = 48'hbc802288a011;
assign testcases[182] = 48'haa801188a001;
assign testcases[183] = 48'hb9700088a000;
assign testcases[184] = 48'hb9700088a000;
assign testcases[185] = 48'hb97000889000;
assign testcases[186] = 48'hb97000889000;
assign testcases[187] = 48'hb97000889000;
assign testcases[188] = 48'hb97000889000;
assign testcases[189] = 48'hb97000889000;
assign testcases[190] = 48'hb97000899000;
assign testcases[191] = 48'hb97000889000;
assign testcases[192] = 48'hd532456b2011;
assign testcases[193] = 48'hb970017a4102;
assign testcases[194] = 48'hb970007a6002;
assign testcases[195] = 48'hb97000898001;
assign testcases[196] = 48'hb97000889000;
assign testcases[197] = 48'hb9700088a000;
assign testcases[198] = 48'hb97000889000;
assign testcases[199] = 48'hb97000889000;
assign testcases[200] = 48'hb97000889000;
assign testcases[201] = 48'hb97000889000;
assign testcases[202] = 48'hb97000889000;
assign testcases[203] = 48'hb9621187f012;
assign testcases[204] = 48'hb9710087d002;
assign testcases[205] = 48'ha9700088b001;
assign testcases[206] = 48'hb97000889000;
assign testcases[207] = 48'hb97000889000;
assign testcases[208] = 48'hb97000899000;
assign testcases[209] = 48'hb97000899000;
assign testcases[210] = 48'hb97000889000;
assign testcases[211] = 48'hb97000889000;
assign testcases[212] = 48'hb97000889000;
assign testcases[213] = 48'hb97000889000;
assign testcases[214] = 48'hb9711197d112;
assign testcases[215] = 48'hb9700087b001;
assign testcases[216] = 48'hb97000889000;
assign testcases[217] = 48'hb97000889000;
assign testcases[218] = 48'hb97000899000;
assign testcases[219] = 48'hb97000889000;
assign testcases[220] = 48'hb97000889000;
assign testcases[221] = 48'hb97000899000;
assign testcases[222] = 48'hb97000889000;
assign testcases[223] = 48'hb97000889000;
assign testcases[224] = 48'hb97000889000;
assign testcases[225] = 48'hb97000889000;
assign testcases[226] = 48'hb97000889000;
assign testcases[227] = 48'hb786765c8555;
assign testcases[228] = 48'ha97786699666;
assign testcases[229] = 48'hb97886889566;
assign testcases[230] = 48'hb9767688a556;
assign testcases[231] = 48'hba758588a455;
assign testcases[232] = 48'hb97686889446;
assign testcases[233] = 48'hc87686899546;
assign testcases[234] = 48'ha97676899555;
assign testcases[235] = 48'hb98676889556;
assign testcases[236] = 48'hc97686889556;
assign testcases[237] = 48'ha96786889556;
assign testcases[238] = 48'haa7685889556;
assign testcases[239] = 48'hc97676899546;
assign testcases[240] = 48'hc97576889546;
assign testcases[241] = 48'hb97575899545;
assign testcases[242] = 48'hc977865b8667;
assign testcases[243] = 48'hb97887699667;
assign testcases[244] = 48'hb97797799677;
assign testcases[245] = 48'hb9769688a666;
assign testcases[246] = 48'haa767688a556;
assign testcases[247] = 48'hc97786889556;
assign testcases[248] = 48'hb97786799656;
assign testcases[249] = 48'hb97786889656;
assign testcases[250] = 48'hc977a7889566;
assign testcases[251] = 48'ha97797889566;
assign testcases[252] = 48'hba7676889466;
assign testcases[253] = 48'hc97676899566;
assign testcases[254] = 48'hb97676899566;
assign testcases[255] = 48'hb97665889455;
assign testcases[256] = 48'hc96c9a899559;
assign testcases[257] = 48'h998c99889568;
assign testcases[258] = 48'hb97ba75b8867;
assign testcases[259] = 48'hb97bb85b8879;
assign testcases[260] = 48'hb97cb879887a;
assign testcases[261] = 48'hca6aa6799778;
assign testcases[262] = 48'hb87bc8a6b788;
assign testcases[263] = 48'hb86cc8b6b788;
assign testcases[264] = 48'hb88ea83e8657;
assign testcases[265] = 48'hb98dc83d7868;
assign testcases[266] = 48'hba6dd93c7868;
assign testcases[267] = 48'hb97dc9889788;
assign testcases[268] = 48'hb96db9799988;
assign testcases[269] = 48'hb87ec9899b88;
assign testcases[270] = 48'ha98dc8c5a878;
assign testcases[271] = 48'ha87ca84d8779;
assign testcases[272] = 48'hd98c985b8689;
assign testcases[273] = 48'hb96ca93d7999;
assign testcases[274] = 48'h987caa699b88;
assign testcases[275] = 48'ha98ca87a9977;
assign testcases[276] = 48'hd97dc8899b88;
assign testcases[277] = 48'hba7dc8c5b779;
assign testcases[278] = 48'hb97db7a7b769;
assign testcases[279] = 48'ha469a84d9457;
assign testcases[280] = 48'hc879a86b8466;
assign testcases[281] = 48'hba7898b58877;
assign testcases[282] = 48'hb97898b59978;
assign testcases[283] = 48'hb86898799457;
assign testcases[284] = 48'hb97788979557;
assign testcases[285] = 48'hb977897aa666;
assign testcases[286] = 48'haa78875d9366;
assign testcases[287] = 48'ha848995b8556;
assign testcases[288] = 48'hb879a8799557;
assign testcases[289] = 48'hc97999a59757;
assign testcases[290] = 48'hb97898b59667;
assign testcases[291] = 48'hb889a8889467;
assign testcases[292] = 48'hba78a8979768;
assign testcases[293] = 48'haa6898799877;
assign testcases[294] = 48'haa79975b9367;
assign testcases[295] = 48'hc849995c8566;
assign testcases[296] = 48'hc97998888667;
assign testcases[297] = 48'hb988a8a69567;
assign testcases[298] = 48'hba79a8999676;
assign testcases[299] = 48'hba7898979676;
assign testcases[300] = 48'hb9788788a867;
assign testcases[301] = 48'ha988874da456;
assign testcases[302] = 48'haad147aaa233;
assign testcases[303] = 48'hb7612488a413;
assign testcases[304] = 48'hb96022789211;
assign testcases[305] = 48'hba8002789111;
assign testcases[306] = 48'hba8012789211;
assign testcases[307] = 48'hb97011889312;
assign testcases[308] = 48'hb97011899112;
assign testcases[309] = 48'hba7011889111;
assign testcases[310] = 48'hb97000889000;
assign testcases[311] = 48'hb97000889000;
assign testcases[312] = 48'hb97000889000;
assign testcases[313] = 48'hb97000889000;
assign testcases[314] = 48'hb97000889100;
assign testcases[315] = 48'hb97000889000;
assign testcases[316] = 48'hb97001889100;
assign testcases[317] = 48'hb97001799301;
assign testcases[318] = 48'hcc7142888101;
assign testcases[319] = 48'hb96001889001;
assign testcases[320] = 48'hb9700088a000;
assign testcases[321] = 48'hb9700089a000;
assign testcases[322] = 48'hb97000899001;
assign testcases[323] = 48'hb97010889000;
assign testcases[324] = 48'hb97010889101;
assign testcases[325] = 48'hb97010889101;
assign testcases[326] = 48'hb97010889000;
assign testcases[327] = 48'hb97000889000;
assign testcases[328] = 48'hb97000889101;
assign testcases[329] = 48'hb95013789411;
assign testcases[330] = 48'hab713188b001;
assign testcases[331] = 48'hb9700088b001;
assign testcases[332] = 48'hb9700088a000;
assign testcases[333] = 48'hb9700088a000;
assign testcases[334] = 48'hb97000889000;
assign testcases[335] = 48'hb97000889000;
assign testcases[336] = 48'hb97000889000;
assign testcases[337] = 48'hb97000889000;
assign testcases[338] = 48'hb97000899000;
assign testcases[339] = 48'hb97000889000;
assign testcases[340] = 48'hb97000889000;
assign testcases[341] = 48'hb9700088a001;
assign testcases[342] = 48'hba7011686101;
assign testcases[343] = 48'hba7000788101;
assign testcases[344] = 48'hb97010789011;
assign testcases[345] = 48'hb9701088a001;
assign testcases[346] = 48'hb9701088a000;
assign testcases[347] = 48'hb97000889000;
assign testcases[348] = 48'hb97000889000;
assign testcases[349] = 48'hb97000899000;
assign testcases[350] = 48'hb97010899001;
assign testcases[351] = 48'hba7010889001;
assign testcases[352] = 48'hb97010889000;
assign testcases[353] = 48'hb9701088a011;
assign testcases[354] = 48'h8a743297f112;
assign testcases[355] = 48'hb9711187c111;
assign testcases[356] = 48'ha9700088b001;
assign testcases[357] = 48'hb9700088a000;
assign testcases[358] = 48'hb97000889000;
assign testcases[359] = 48'hb97000889000;
assign testcases[360] = 48'hb97000889000;
assign testcases[361] = 48'hb97000899000;
assign testcases[362] = 48'hb97000889000;
assign testcases[363] = 48'hb97000889000;
assign testcases[364] = 48'hb97000889000;
assign testcases[365] = 48'hb97000889000;
assign testcases[366] = 48'hb97000889000;
assign testcases[367] = 48'hb97000889000;
assign testcases[368] = 48'hb97000899000;
assign testcases[369] = 48'hb97000889011;
assign testcases[370] = 48'hc9623297e212;
assign testcases[371] = 48'hca612297c212;
assign testcases[372] = 48'hb9700188a001;
assign testcases[373] = 48'hb97000889000;
assign testcases[374] = 48'hb97000889000;
assign testcases[375] = 48'hb97000899000;
assign testcases[376] = 48'hb97000899000;
assign testcases[377] = 48'hb97000889000;
assign testcases[378] = 48'hb97000889000;
assign testcases[379] = 48'hb97000889000;
assign testcases[380] = 48'hb97000889000;
assign testcases[381] = 48'hb97000889000;
assign testcases[382] = 48'hb97000889000;
assign testcases[383] = 48'hb97000889000;
assign testcases[384] = 48'hbb7565698434;
assign testcases[385] = 48'hb97674799544;
assign testcases[386] = 48'hb9766579a544;
assign testcases[387] = 48'hb97665889443;
assign testcases[388] = 48'hb97674889543;
assign testcases[389] = 48'hca7674899544;
assign testcases[390] = 48'hb97675899545;
assign testcases[391] = 48'hb87675889544;
assign testcases[392] = 48'hb96685889544;
assign testcases[393] = 48'hb97574889534;
assign testcases[394] = 48'hc97674899434;
assign testcases[395] = 48'hba866589a334;
assign testcases[396] = 48'hb97666799433;
assign testcases[397] = 48'hb87575889543;
assign testcases[398] = 48'hba7565889544;
assign testcases[399] = 48'hca7574889534;
assign testcases[400] = 48'hb86676b89545;
assign testcases[401] = 48'hb97675989535;
assign testcases[402] = 48'hba7684799535;
assign testcases[403] = 48'hb9767579a544;
assign testcases[404] = 48'hb87675889535;
assign testcases[405] = 48'hba7685889645;
assign testcases[406] = 48'hca7685889644;
assign testcases[407] = 48'hb97685799545;
assign testcases[408] = 48'hb87675889644;
assign testcases[409] = 48'hb97685889544;
assign testcases[410] = 48'hca7685889544;
assign testcases[411] = 48'hb97675799544;
assign testcases[412] = 48'hb97665899534;
assign testcases[413] = 48'hb97675889444;
assign testcases[414] = 48'hba7685889544;
assign testcases[415] = 48'hca8a55889535;
assign testcases[416] = 48'haa7955789535;
assign testcases[417] = 48'hc97a66498835;
assign testcases[418] = 48'haa8b54b8a435;
assign testcases[419] = 48'hb97c54a8a435;
assign testcases[420] = 48'haa88455a8435;
assign testcases[421] = 48'hba8945799435;
assign testcases[422] = 48'hc97955699435;
assign testcases[423] = 48'hc87875498835;
assign testcases[424] = 48'hb97875689a36;
assign testcases[425] = 48'h998856899735;
assign testcases[426] = 48'ha97867799846;
assign testcases[427] = 48'ha96956a8a546;
assign testcases[428] = 48'hb97b55a7a435;
assign testcases[429] = 48'he96c6669aa35;
assign testcases[430] = 48'hca8b565a8545;
assign testcases[431] = 48'haa8b55689535;
assign testcases[432] = 48'ha97a65498736;
assign testcases[433] = 48'ha87965698936;
assign testcases[434] = 48'hba7a56799845;
assign testcases[435] = 48'hb97966799945;
assign testcases[436] = 48'hc97b74b6a636;
assign testcases[437] = 48'hca6c65b8b536;
assign testcases[438] = 48'hc75887878348;
assign testcases[439] = 48'haa7866789448;
assign testcases[440] = 48'h998866989448;
assign testcases[441] = 48'hb98877b8b546;
assign testcases[442] = 48'hb9677799a647;
assign testcases[443] = 48'hc96875698449;
assign testcases[444] = 48'hb97776979749;
assign testcases[445] = 48'ha97776979649;
assign testcases[446] = 48'hc878766a9449;
assign testcases[447] = 48'hc978766aa447;
assign testcases[448] = 48'haa77666aa547;
assign testcases[449] = 48'ha6797698a548;
assign testcases[450] = 48'hb97966889547;
assign testcases[451] = 48'hc98877a8a656;
assign testcases[452] = 48'hc97886b7b656;
assign testcases[453] = 48'hb96876889757;
assign testcases[454] = 48'hb9798798a658;
assign testcases[455] = 48'hb97987899658;
assign testcases[456] = 48'hb879875a8558;
assign testcases[457] = 48'hb97986699658;
assign testcases[458] = 48'hc66a97b9a658;
assign testcases[459] = 48'hc88a76999657;
assign testcases[460] = 48'hb97877b6a658;
assign testcases[461] = 48'hb97987a79858;
assign testcases[462] = 48'hb97986799758;
assign testcases[463] = 48'hb9898897a758;
assign testcases[464] = 48'hb96978699857;
assign testcases[465] = 48'hb969774b9657;
assign testcases[466] = 48'hcfe3758f4146;
assign testcases[467] = 48'ha991268b9123;
assign testcases[468] = 48'hb86011899212;
assign testcases[469] = 48'hb96012789112;
assign testcases[470] = 48'hb9702188a102;
assign testcases[471] = 48'hb9701188a101;
assign testcases[472] = 48'hb97000889101;
assign testcases[473] = 48'hb97010789101;
assign testcases[474] = 48'hb97010899101;
assign testcases[475] = 48'hb97011899101;
assign testcases[476] = 48'hb98011899101;
assign testcases[477] = 48'hb97011889101;
assign testcases[478] = 48'hb97011889101;
assign testcases[479] = 48'hb97001889000;
assign testcases[480] = 48'hb97001889000;
assign testcases[481] = 48'hb8702188a111;
assign testcases[482] = 48'hde8172887212;
assign testcases[483] = 48'hb87021888101;
assign testcases[484] = 48'hb97011789101;
assign testcases[485] = 48'hb97010889201;
assign testcases[486] = 48'hba7020899201;
assign testcases[487] = 48'hba702178a101;
assign testcases[488] = 48'hb8701088a101;
assign testcases[489] = 48'hb97011889101;
assign testcases[490] = 48'hba6010889001;
assign testcases[491] = 48'hb9701189a001;
assign testcases[492] = 48'hb88000899000;
assign testcases[493] = 48'hb97011889101;
assign testcases[494] = 48'h8d719188d011;
assign testcases[495] = 48'hb8701088c001;
assign testcases[496] = 48'hb9700088b001;
assign testcases[497] = 48'hb9700088a001;
assign testcases[498] = 48'hb97000889000;
assign testcases[499] = 48'hb97010899001;
assign testcases[500] = 48'hb97011899001;
assign testcases[501] = 48'hb97010889011;
assign testcases[502] = 48'hb97011889011;
assign testcases[503] = 48'hb96000889010;
assign testcases[504] = 48'hb97000889000;
assign testcases[505] = 48'hb97000899000;
assign testcases[506] = 48'hb97000889000;
assign testcases[507] = 48'hb97000889000;
assign testcases[508] = 48'hbda159575315;
assign testcases[509] = 48'hb85011678112;
assign testcases[510] = 48'hb87010789101;
assign testcases[511] = 48'hb97010889101;
assign testcases[512] = 48'hb97010889001;
assign testcases[513] = 48'hba7010899001;
assign testcases[514] = 48'hb97011899111;
assign testcases[515] = 48'hba8011899111;
assign testcases[516] = 48'hbb7011889011;
assign testcases[517] = 48'hb8713288a023;
assign testcases[518] = 48'hb8813289a023;
assign testcases[519] = 48'hb97012889121;
assign testcases[520] = 48'h4b864299f112;
assign testcases[521] = 48'hc9711099d111;
assign testcases[522] = 48'hb9700088b001;
assign testcases[523] = 48'hb9701088a001;
assign testcases[524] = 48'hb97011889111;
assign testcases[525] = 48'hb97011889001;
assign testcases[526] = 48'hb97000889000;
assign testcases[527] = 48'hb97000889000;
assign testcases[528] = 48'hb97000899000;
assign testcases[529] = 48'hb97000889000;
assign testcases[530] = 48'hb97000889000;
assign testcases[531] = 48'hb97010899000;
assign testcases[532] = 48'h89843298f111;
assign testcases[533] = 48'hc9711188d112;
assign testcases[534] = 48'hb9700088b001;
assign testcases[535] = 48'hb9700088a001;
assign testcases[536] = 48'hb97000889000;
assign testcases[537] = 48'hb97000889000;
assign testcases[538] = 48'hb97000889000;
assign testcases[539] = 48'hb97000889000;
assign testcases[540] = 48'hb97000899000;
assign testcases[541] = 48'hb97000889000;
assign testcases[542] = 48'hb97000889000;
assign testcases[543] = 48'hb97000899000;
assign testcases[544] = 48'hb96674888434;
assign testcases[545] = 48'hba767479a533;
assign testcases[546] = 48'hb87674799543;
assign testcases[547] = 48'hb97684889543;
assign testcases[548] = 48'hba7784889643;
assign testcases[549] = 48'hb97684799644;
assign testcases[550] = 48'hb97684889643;
assign testcases[551] = 48'hba7684889643;
assign testcases[552] = 48'hc97684889633;
assign testcases[553] = 48'hb88674799543;
assign testcases[554] = 48'hb97684899543;
assign testcases[555] = 48'hb97684889543;
assign testcases[556] = 48'hb97784889543;
assign testcases[557] = 48'hb97774799543;
assign testcases[558] = 48'hba6574298e44;
assign testcases[559] = 48'hb87684b8a544;
assign testcases[560] = 48'hba677498a643;
assign testcases[561] = 48'hb97784799633;
assign testcases[562] = 48'hb97794889634;
assign testcases[563] = 48'hb97794889644;
assign testcases[564] = 48'hb977847a9644;
assign testcases[565] = 48'ha97784899643;
assign testcases[566] = 48'hb97694889533;
assign testcases[567] = 48'hb96784889643;
assign testcases[568] = 48'hb97784799743;
assign testcases[569] = 48'ha98784889743;
assign testcases[570] = 48'hb97694889643;
assign testcases[571] = 48'hc96693899643;
assign testcases[572] = 48'hba8674799643;
assign testcases[573] = 48'hc97c66788535;
assign testcases[574] = 48'hca8c66789534;
assign testcases[575] = 48'hc87b86488736;
assign testcases[576] = 48'ha97b86789947;
assign testcases[577] = 48'haa7a6679a845;
assign testcases[578] = 48'ha86b76889935;
assign testcases[579] = 48'ha97d66b8a535;
assign testcases[580] = 48'hca6e6599a635;
assign testcases[581] = 48'hba7d66698636;
assign testcases[582] = 48'hba6c655a8535;
assign testcases[583] = 48'hb87b76497946;
assign testcases[584] = 48'hd98c86688a37;
assign testcases[585] = 48'hc97c86789936;
assign testcases[586] = 48'h987d8597a936;
assign testcases[587] = 48'haa6f76b7b635;
assign testcases[588] = 48'hca7e66598535;
assign testcases[589] = 48'hba7d864a8645;
assign testcases[590] = 48'hc87c87498a47;
assign testcases[591] = 48'hb97c76688a47;
assign testcases[592] = 48'h9a8c76789835;
assign testcases[593] = 48'hc97d77a7a838;
assign testcases[594] = 48'hb95d96b8b748;
assign testcases[595] = 48'ha66a88b89567;
assign testcases[596] = 48'hb98978a89566;
assign testcases[597] = 48'hca8978b6a666;
assign testcases[598] = 48'hb97978989766;
assign testcases[599] = 48'hb87987789667;
assign testcases[600] = 48'hb87986979757;
assign testcases[601] = 48'ha96977698866;
assign testcases[602] = 48'ha969774a9666;
assign testcases[603] = 48'hb67a87a8a657;
assign testcases[604] = 48'hc97a87989566;
assign testcases[605] = 48'hc97986b7a567;
assign testcases[606] = 48'hb97987a89757;
assign testcases[607] = 48'ha98987889566;
assign testcases[608] = 48'hb9788798a666;
assign testcases[609] = 48'haa69876b9755;
assign testcases[610] = 48'haa79875a9556;
assign testcases[611] = 48'hb46a97c8a756;
assign testcases[612] = 48'ha97a87b89755;
assign testcases[613] = 48'haa7987c69668;
assign testcases[614] = 48'hb98987a89868;
assign testcases[615] = 48'hca887889a756;
assign testcases[616] = 48'hb87977889665;
assign testcases[617] = 48'ha87977499565;
assign testcases[618] = 48'ha96977698766;
assign testcases[619] = 48'hba811289a121;
assign testcases[620] = 48'hb9700188a101;
assign testcases[621] = 48'hb97001899000;
assign testcases[622] = 48'hb97001889000;
assign testcases[623] = 48'hb97001889000;
assign testcases[624] = 48'hb97000889000;
assign testcases[625] = 48'hb97000889000;
assign testcases[626] = 48'hb97000899000;
assign testcases[627] = 48'hb97000889000;
assign testcases[628] = 48'hb97000889000;
assign testcases[629] = 48'hb98003889100;
assign testcases[630] = 48'hb97001889100;
assign testcases[631] = 48'hb97000889000;
assign testcases[632] = 48'hb97000889000;
assign testcases[633] = 48'hb97000889000;
assign testcases[634] = 48'hb97000889000;
assign testcases[635] = 48'hb97000889000;
assign testcases[636] = 48'hb97010799301;
assign testcases[637] = 48'hb86111889422;
assign testcases[638] = 48'hb96112889222;
assign testcases[639] = 48'hba8011899111;
assign testcases[640] = 48'hba8012899111;
assign testcases[641] = 48'ha9812288a111;
assign testcases[642] = 48'hb9700188a000;
assign testcases[643] = 48'hb9700088a000;
assign testcases[644] = 48'hb97000889000;
assign testcases[645] = 48'hb97000899000;
assign testcases[646] = 48'hb97000889000;
assign testcases[647] = 48'hb97000889000;
assign testcases[648] = 48'hb97000889000;
assign testcases[649] = 48'hb97000889000;
assign testcases[650] = 48'hb97000889000;
assign testcases[651] = 48'hb97000889000;
assign testcases[652] = 48'hb981126e7111;
assign testcases[653] = 48'hb970017b9111;
assign testcases[654] = 48'hb97001799010;
assign testcases[655] = 48'hb97000889000;
assign testcases[656] = 48'hb97001889000;
assign testcases[657] = 48'hb97011889010;
assign testcases[658] = 48'hb97011889000;
assign testcases[659] = 48'hba7011889001;
assign testcases[660] = 48'hb97011899010;
assign testcases[661] = 48'hb97011889010;
assign testcases[662] = 48'hb97011889010;
assign testcases[663] = 48'hb97001899000;
assign testcases[664] = 48'hb97001889000;
assign testcases[665] = 48'hb97000889000;
assign testcases[666] = 48'h29883482c221;
assign testcases[667] = 48'hc9711284b131;
assign testcases[668] = 48'hb9711286a121;
assign testcases[669] = 48'ha97101889111;
assign testcases[670] = 48'ha97101899010;
assign testcases[671] = 48'ha97100889000;
assign testcases[672] = 48'hb97000889000;
assign testcases[673] = 48'hb97000889010;
assign testcases[674] = 48'hb97000889010;
assign testcases[675] = 48'hb97000889000;
assign testcases[676] = 48'hb97000889000;
assign testcases[677] = 48'hb97000889000;
assign testcases[678] = 48'h97713193c212;
assign testcases[679] = 48'ha8711195b111;
assign testcases[680] = 48'hb9700087a011;
assign testcases[681] = 48'hb97010889010;
assign testcases[682] = 48'hb97000899000;
assign testcases[683] = 48'hc97111889110;
assign testcases[684] = 48'hb97111899111;
assign testcases[685] = 48'hb97010899111;
assign testcases[686] = 48'hb97111899110;
assign testcases[687] = 48'ha97111899110;
assign testcases[688] = 48'hb97100889010;
assign testcases[689] = 48'hb97000889000;
assign testcases[690] = 48'hb8687a8aa558;
assign testcases[691] = 48'hb9887a899658;
assign testcases[692] = 48'hba787a988668;
assign testcases[693] = 48'hb9797a889659;
assign testcases[694] = 48'hb9797a79a659;
assign testcases[695] = 48'hb9787b899758;
assign testcases[696] = 48'hba887a889758;
assign testcases[697] = 48'hb97759889547;
assign testcases[698] = 48'hb9765a98a546;
assign testcases[699] = 48'hb9766a789646;
assign testcases[700] = 48'haa7669789546;
assign testcases[701] = 48'hc9766a899557;
assign testcases[702] = 48'hb9776a889547;
assign testcases[703] = 48'ha8686b3ba656;
assign testcases[704] = 48'hb9786a49a647;
assign testcases[705] = 48'hb96879799648;
assign testcases[706] = 48'hba7769888548;
assign testcases[707] = 48'hb9786a889558;
assign testcases[708] = 48'hb8787a89a658;
assign testcases[709] = 48'hb9787a899768;
assign testcases[710] = 48'hba788a989758;
assign testcases[711] = 48'hba897a889658;
assign testcases[712] = 48'hb9887978a558;
assign testcases[713] = 48'hb87869799548;
assign testcases[714] = 48'ha97779899658;
assign testcases[715] = 48'hba7779989447;
assign testcases[716] = 48'hc99b66899456;
assign testcases[717] = 48'hc97d66689656;
assign testcases[718] = 48'hc98d56999957;
assign testcases[719] = 48'hd95c57699868;
assign testcases[720] = 48'h9a8b57999758;
assign testcases[721] = 48'hb98c67b8a556;
assign testcases[722] = 48'hd86d67889667;
assign testcases[723] = 48'ha976660bc557;
assign testcases[724] = 48'hb8666649a548;
assign testcases[725] = 48'hc95666688448;
assign testcases[726] = 48'ha86456798438;
assign testcases[727] = 48'hba7667a8a959;
assign testcases[728] = 48'ha8665788984a;
assign testcases[729] = 48'hc9866798974a;
assign testcases[730] = 48'hca865659a54a;
assign testcases[731] = 48'hb9765649b549;
assign testcases[732] = 48'ha96666a98c59;
assign testcases[733] = 48'haa8c673aa658;
assign testcases[734] = 48'hb97c6658b567;
assign testcases[735] = 48'hbaaca96ab689;
assign testcases[736] = 48'hb88daa699989;
assign testcases[737] = 48'hc97e8a888a8a;
assign testcases[738] = 48'haa7e68b8a578;
assign testcases[739] = 48'hb757663aa64a;
assign testcases[740] = 48'hb767566aa74b;
assign testcases[741] = 48'ha97678a9885d;
assign testcases[742] = 48'hba777898976c;
assign testcases[743] = 48'hba8656899659;
assign testcases[744] = 48'hb97656a8955a;
assign testcases[745] = 48'hc8676668b75b;
assign testcases[746] = 48'hc8776659a65a;
assign testcases[747] = 48'haa9d674aa777;
assign testcases[748] = 48'hd98e6748a766;
assign testcases[749] = 48'hc86e78399666;
assign testcases[750] = 48'ha96f8b788987;
assign testcases[751] = 48'hb85fac79aa88;
assign testcases[752] = 48'hba9daa8a9978;
assign testcases[753] = 48'habae78c79568;
assign testcases[754] = 48'hb87f67b7a587;
assign testcases[755] = 48'hb856672ba64b;
assign testcases[756] = 48'ha965663a864b;
assign testcases[757] = 48'hb9767798695b;
assign testcases[758] = 48'hca7777a8985c;
assign testcases[759] = 48'hb9777699a65c;
assign testcases[760] = 48'ha8767798a55c;
assign testcases[761] = 48'hb9767768b56b;
assign testcases[762] = 48'hb975665ab55a;
assign testcases[763] = 48'hc7a24479b434;
assign testcases[764] = 48'hc78124889212;
assign testcases[765] = 48'hb86011889111;
assign testcases[766] = 48'hb97011889100;
assign testcases[767] = 48'hb98001889100;
assign testcases[768] = 48'hb97000889000;
assign testcases[769] = 48'hb97000889000;
assign testcases[770] = 48'hb97000889100;
assign testcases[771] = 48'hb97000889100;
assign testcases[772] = 48'hb97000889000;
assign testcases[773] = 48'hb97000889000;
assign testcases[774] = 48'hb9a1248cc233;
assign testcases[775] = 48'hb970128ab112;
assign testcases[776] = 48'hb9701189a011;
assign testcases[777] = 48'hb97000889000;
assign testcases[778] = 48'hb97000889000;
assign testcases[779] = 48'hb97001889111;
assign testcases[780] = 48'hb97101889111;
assign testcases[781] = 48'hb97001889011;
assign testcases[782] = 48'hb97000889000;
assign testcases[783] = 48'hb97000889000;
assign testcases[784] = 48'hb97000889000;
assign testcases[785] = 48'hb97000899000;
assign testcases[786] = 48'hb99137877111;
assign testcases[787] = 48'hba6012878001;
assign testcases[788] = 48'hb97000889001;
assign testcases[789] = 48'ha6b1478aa122;
assign testcases[790] = 48'ha7926a889144;
assign testcases[791] = 48'h87a47d8aa166;
assign testcases[792] = 48'h34f36a8bb245;
assign testcases[793] = 48'h77b337868212;
assign testcases[794] = 48'hb97111868011;
assign testcases[795] = 48'hb97011878011;
assign testcases[796] = 48'hb97111889111;
assign testcases[797] = 48'hb97111899011;
assign testcases[798] = 48'ha971226fb121;
assign testcases[799] = 48'hb970117da111;
assign testcases[800] = 48'hb970117aa111;
assign testcases[801] = 48'hb97001899001;
assign testcases[802] = 48'hb97000889000;
assign testcases[803] = 48'hb97000889000;
assign testcases[804] = 48'hb97001889000;
assign testcases[805] = 48'hb97000889000;
assign testcases[806] = 48'hb98112899010;
assign testcases[807] = 48'hb98112889121;
assign testcases[808] = 48'hb97012889111;
assign testcases[809] = 48'hb97011899001;
assign testcases[810] = 48'hb97000899000;
assign testcases[811] = 48'hc97101848111;
assign testcases[812] = 48'hb97000879010;
assign testcases[813] = 48'hb97000889000;
assign testcases[814] = 48'hb97000899100;
assign testcases[815] = 48'hb97011899111;
assign testcases[816] = 48'hb9711189a211;
assign testcases[817] = 48'ha97111899211;
assign testcases[818] = 48'hb97011889110;
assign testcases[819] = 48'hb97011889000;
assign testcases[820] = 48'hb97000889000;
assign testcases[821] = 48'hb97000889000;
assign testcases[822] = 48'hc96101928120;
assign testcases[823] = 48'hb97000868110;
assign testcases[824] = 48'hb97000889010;
assign testcases[825] = 48'hb97000899000;
assign testcases[826] = 48'hb97111899110;
assign testcases[827] = 48'haa8111899110;
assign testcases[828] = 48'hba7111889000;
assign testcases[829] = 48'hb97010889000;
assign testcases[830] = 48'hb97011889111;
assign testcases[831] = 48'hb97011889111;
assign testcases[832] = 48'hb97000899000;
assign testcases[833] = 48'hb97000889000;
assign testcases[834] = 48'hb97010889011;
assign testcases[835] = 48'hc97111889111;
assign testcases[836] = 48'hb87111789111;
assign testcases[837] = 48'hba796a3ad578;
assign testcases[838] = 48'hb9796a58a779;
assign testcases[839] = 48'hb9696a78a789;
assign testcases[840] = 48'hb97a7b89a789;
assign testcases[841] = 48'hb9897b99977a;
assign testcases[842] = 48'hba787a988679;
assign testcases[843] = 48'hb9797978a779;
assign testcases[844] = 48'hb9697a78a678;
assign testcases[845] = 48'hb9797c999589;
assign testcases[846] = 48'hb9897c89868a;
assign testcases[847] = 48'hba796b889579;
assign testcases[848] = 48'hb9796a78a568;
assign testcases[849] = 48'hc9796979a679;
assign testcases[850] = 48'hc9796a38e378;
assign testcases[851] = 48'hb9796b59c578;
assign testcases[852] = 48'hb9895b799568;
assign testcases[853] = 48'hb9795a989578;
assign testcases[854] = 48'hb9795987a568;
assign testcases[855] = 48'hb9796a79a578;
assign testcases[856] = 48'ha97a6a899689;
assign testcases[857] = 48'hb9796a988578;
assign testcases[858] = 48'hba796a88a678;
assign testcases[859] = 48'hb9796b78a578;
assign testcases[860] = 48'hb9696b899578;
assign testcases[861] = 48'hb9796b898588;
assign testcases[862] = 48'hc9796b889689;
assign testcases[863] = 48'hc97d5c78a677;
assign testcases[864] = 48'hc96d5c58b677;
assign testcases[865] = 48'h988c6c49b577;
assign testcases[866] = 48'hc98e7c899688;
assign testcases[867] = 48'hca7d6d7897a9;
assign testcases[868] = 48'ha97c6e8898aa;
assign testcases[869] = 48'hca7e7dc8748b;
assign testcases[870] = 48'hc87e5fb97599;
assign testcases[871] = 48'hb87e5e69a788;
assign testcases[872] = 48'ha96e6f49b688;
assign testcases[873] = 48'hba7e6f799688;
assign testcases[874] = 48'ha99d5d69a788;
assign testcases[875] = 48'hd97d5d89998a;
assign testcases[876] = 48'hc97e6cb8757a;
assign testcases[877] = 48'hac676a49cb8b;
assign testcases[878] = 48'ha9775919d788;
assign testcases[879] = 48'hb8786a8a7a9a;
assign testcases[880] = 48'hba886aa9889a;
assign testcases[881] = 48'hb9885a88b888;
assign testcases[882] = 48'hb86869979798;
assign testcases[883] = 48'hba675867b788;
assign testcases[884] = 48'hb9775858b778;
assign testcases[885] = 48'h9c686939d789;
assign testcases[886] = 48'ha9794939d799;
assign testcases[887] = 48'hb8785a8979aa;
assign testcases[888] = 48'ha9775aa9899a;
assign testcases[889] = 48'ha9775998a998;
assign testcases[890] = 48'hc8685a9997a9;
assign testcases[891] = 48'hda795a68b898;
assign testcases[892] = 48'haa794b48c896;
assign testcases[893] = 48'ha9884a5ab897;
assign testcases[894] = 48'hc9786aa9789b;
assign testcases[895] = 48'hb97769a9889c;
assign testcases[896] = 48'ha97859989988;
assign testcases[897] = 48'hc8695b988798;
assign testcases[898] = 48'hca685b68b898;
assign testcases[899] = 48'hb9784a48c796;
assign testcases[900] = 48'hd88d5c47c588;
assign testcases[901] = 48'hc96d6d47b588;
assign testcases[902] = 48'ha97c6e38b578;
assign testcases[903] = 48'hc97d6e899779;
assign testcases[904] = 48'hd96e7f78a799;
assign testcases[905] = 48'h998e7f8998a9;
assign testcases[906] = 48'hb98f5eb97588;
assign testcases[907] = 48'hba802288a311;
assign testcases[908] = 48'hb9712178a212;
assign testcases[909] = 48'hb9712178a111;
assign testcases[910] = 48'hb9701088a101;
assign testcases[911] = 48'hb97010889100;
assign testcases[912] = 48'hb97010899100;
assign testcases[913] = 48'hb97000889000;
assign testcases[914] = 48'hb97000889000;
assign testcases[915] = 48'hb97000889100;
assign testcases[916] = 48'hb97000889000;
assign testcases[917] = 48'hb97000889000;
assign testcases[918] = 48'hb97000889000;
assign testcases[919] = 48'hb96111898111;
assign testcases[920] = 48'hb97000899000;
assign testcases[921] = 48'hb97000899000;
assign testcases[922] = 48'hb97000889000;
assign testcases[923] = 48'hb97000889000;
assign testcases[924] = 48'hb97000889000;
assign testcases[925] = 48'hb97000889000;
assign testcases[926] = 48'hb97000889000;
assign testcases[927] = 48'hb97000889000;
assign testcases[928] = 48'hb97000899000;
assign testcases[929] = 48'hb98011899111;
assign testcases[930] = 48'h9c827177d001;
assign testcases[931] = 48'hb8702088c001;
assign testcases[932] = 48'hb9700088b001;
assign testcases[933] = 48'hb9700088a000;
assign testcases[934] = 48'hb97000889000;
assign testcases[935] = 48'hb97000889000;
assign testcases[936] = 48'hb97000889000;
assign testcases[937] = 48'hb97000889000;
assign testcases[938] = 48'hb97000889000;
assign testcases[939] = 48'hb97000889000;
assign testcases[940] = 48'hb97000889000;
assign testcases[941] = 48'hb97000889000;
assign testcases[942] = 48'h9e7152773113;
assign testcases[943] = 48'hb97120786002;
assign testcases[944] = 48'hb97010788001;
assign testcases[945] = 48'hb97000899000;
assign testcases[946] = 48'hb9700089a000;
assign testcases[947] = 48'hb9700088a000;
assign testcases[948] = 48'hb97000889000;
assign testcases[949] = 48'hb97000889000;
assign testcases[950] = 48'hb97000889000;
assign testcases[951] = 48'hb97000889000;
assign testcases[952] = 48'hb97000889000;
assign testcases[953] = 48'hb97000889000;
assign testcases[954] = 48'hf9632288e144;
assign testcases[955] = 48'hb9710089b011;
assign testcases[956] = 48'hb97000899001;
assign testcases[957] = 48'hb97000889000;
assign testcases[958] = 48'hb97000889000;
assign testcases[959] = 48'hb97000889000;
assign testcases[960] = 48'hb97000889000;
assign testcases[961] = 48'hb97000889000;
assign testcases[962] = 48'hb97000889000;
assign testcases[963] = 48'hb97000889000;
assign testcases[964] = 48'hb97000889000;
assign testcases[965] = 48'hb97000889000;
assign testcases[966] = 48'hb97000889000;
assign testcases[967] = 48'hb97000899000;
assign testcases[968] = 48'hb97000889000;
assign testcases[969] = 48'h8004798fc622;
assign testcases[970] = 48'hc871228cb411;
assign testcases[971] = 48'hb970017aa111;
assign testcases[972] = 48'hb9700179a100;
assign testcases[973] = 48'hb97000789000;
assign testcases[974] = 48'hba7010889000;
assign testcases[975] = 48'hb97010889000;
assign testcases[976] = 48'hb87010889000;
assign testcases[977] = 48'hb97000889000;
assign testcases[978] = 48'hb97000889000;
assign testcases[979] = 48'hb97000889000;
assign testcases[980] = 48'hb97000889000;
assign testcases[981] = 48'hb97000889000;
assign testcases[982] = 48'hb97000889000;
assign testcases[983] = 48'hb97000889000;
assign testcases[984] = 48'hb97011889100;
assign testcases[985] = 48'ha97896a79779;
assign testcases[986] = 48'hca899788967a;
assign testcases[987] = 48'hc97a9688977a;
assign testcases[988] = 48'ha9799788a88a;
assign testcases[989] = 48'hba689779a78a;
assign testcases[990] = 48'hc8789779968b;
assign testcases[991] = 48'hb8789789878a;
assign testcases[992] = 48'haa7897799789;
assign testcases[993] = 48'hc9899788968a;
assign testcases[994] = 48'hc9798789978a;
assign testcases[995] = 48'ha9798688a78a;
assign testcases[996] = 48'hb9779688a779;
assign testcases[997] = 48'hca77a6889779;
assign testcases[998] = 48'hc877a7788679;
assign testcases[999] = 48'ha98786a7a779;



Har_bnn1_bnnpar dut (.features(features),.prediction(prediction));

integer i;
initial begin
    features = testcases[0];
    $write("[");//"
    for(i=0;i<TEST_CNT;i=i+1) begin
        features = testcases[i];
        #period
        $write("%d, ",prediction);
    end
    $display("]");
end

endmodule
