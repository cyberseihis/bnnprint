
















module Har_tnn1_tnnpaarter #(

parameter FEAT_CNT = 12,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 5664'h002500650001000300630001000e00610001003b005d00010037005c00010024005b0001001100570001001a00550001002b005400010008005300010015005200010043005100010003004f00010048004e0001003d004c00010001004900010035004200010016003c0001000b002c00010007002b0001002000290001000f00260001000f00220001000000220001001400160001000f00130001002d005000000041004d0000001c004700000032004600000017004500000020004400000011004000000033003f00000026003e00000024003a0000002e00390000001700360000001b003400000021003100000004003000000012002f00000023002e0000001f002d00000028002c00000016002a0000001d00290000000800280000001c00270000000900270000001000250000000500210000001a001f00000015001f0000001c001e00000015001e0000000f001e00000013001b0000000f001a0000001300170000000f00160000000d00130000000800130000000100130000000500100000000100100000000e000f00000008000f00000007000e00000004000e0000000a000d00000004000c00000006000b00000004000b00000007000a00000000000900000004000600000001000300000000000200000016002a00010005001a00010011002300000006000d00000009001b0001000a001800010000001800010002001400010008001100010003000d00010007000c00010005000700010019001d0000000c00190000000f00150000000d00140000000e001200000001000200000011001700010001000c00010003001200000002000900000001000200010004000800010003000a0000000000050000000400080000000b001000010005000d0001000000050001000b000e00000003000900000008000c00010006000700010002000400010006000700000003000a00010000000100010009000b0000 ;
localparam YMAP = 1280'h0000007a0001006f0000006c000000700000007e0001005900010080000000660001007c000000780000006d00000077000100710000007f00010062000100720000007d000000670000006800010056000000790001004a000000580000006a0001006900010060000000730001005e0000006e00000074000000810000005a000000640001004b0001005f0000006b0000007500000038000000760001007b;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 240'b100000010000110000000010001010000000100100000001000000000000000001011001001000000000010110000001001000110000000000010001000000010000101100000110000001000100001000000100000000010001010001010100010000000000010000000011000100100010010001000000 ;
localparam WNNZ = 240'b110010010010110010000110001010000000100101001001101000100000010001011001001100000100010110100001001001110000100000010011000000110000111101100110001001000100001100011110101000010101010101011100011000000001010101010111010100110110010001000000;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
wire [SUM_BITS-1:0] scorarr [CLASS_CNT-1:0];
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;

generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam adsub = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(adsub)
        assign node[nodeloc] = node[op1] - node[op2];
    else
        assign node[nodeloc] = node[op1] + node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] <= 0;
end
endgenerate

function [7:0] zerocnt(input integer k);
    integer i,j;
    reg [HIDDEN_CNT-1:0] neur1;
    begin
        i = 0;
        neur1 = WNNZ[k*HIDDEN_CNT+:HIDDEN_CNT];
        for(j=0;j<HIDDEN_CNT;j=j+1)
            i = i + !(neur1[j]);
        zerocnt = i;
    end
endfunction

function [7:0] minzc(input integer k);
    integer i,j,h;
    begin
        i = HIDDEN_CNT;
        for(j=0;j<CLASS_CNT;j=j+1) begin
            h = zerocnt(j);
            if(h<i)
                i = h;
        end
        minzc = i;
    end
endfunction

localparam MINZC = minzc(0);

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    localparam Wuse = WNNZ[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wuse[j]) begin
            if(Wneur[j])
                tmpscore = tmpscore + hidden[j];
            else 
                tmpscore = tmpscore + hidden_n[j];
        end
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = 2*tmpscore + zerocnt(i) - MINZC;
    /* assign scorarr[i] = 2*tmpscore + zerocnt(i) - MINZC; */
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
