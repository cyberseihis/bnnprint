











module winered_tnn1_tnnzeq #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnnzeq #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(440'b00011100000000110110110000000000000000011001010001000010000100000111001000000101001011010001000100010100000101000010100110001000011010000010001001001011011000010100000010110100001001001011100101000100000101000010100000001001010000010111100100010010001011001000000000001000010000111011101010110010110000000010100000000000100000000010000001111000010111101001000010000000000000010011001100000001011000101010000000000000000010100000001000100100),
  .MASK(440'b11111100100001110110110000001001000010111011011111011011110100010111001011101101101011111101000101011111100101010010101110101100011010001010101111101111111010110101011110111100001011111111100101001111100111001010100001011111110000110111110100110011101011011010111001101000010000111111101110110011111010100110100111001100101100011010000101111110010111111001111010101001001010011111001111111011011010101110000010001100101010110100101011111111),
  .NONZERO_CNT(640'h070702060806070805080605050a0608080607040707070704070806060506080704080805040609),
  .SPARSE_VALS2(71'b11111010010011110001001011010000111010010110011001101111011010010001010),  // Bits of not-zeroes
  .COL_INDICES(568'h2523211e190e0d0c08060400252421201f1d1916140f0e0c0b070302010027222120170c06012321190e0d0c0908040100231d1c0d0b0a0905271e1d1c1a171612110c04030200), // Column of non-zeros
  .ROW_PTRS(56'h473b2921160e00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
