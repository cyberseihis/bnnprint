`timescale 1us/1ns









module tbwinered_tnn1_tnnpar #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


)();
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
reg clk;
reg [FEAT_CNT*FEAT_BITS-1:0] features;
wire [$clog2(CLASS_CNT)-1:0] prediction;
wire [FEAT_CNT*FEAT_BITS-1:0] testcases [TEST_CNT-1:0];
parameter Nsperiod=5000;
localparam period=Nsperiod/500;


assign testcases[0] = 44'h22a92221064;
assign testcases[1] = 44'h33683522085;
assign testcases[2] = 44'h33783322175;
assign testcases[3] = 44'h32593421929;
assign testcases[4] = 44'h22a92221064;
assign testcases[5] = 44'h22a92321064;
assign testcases[6] = 44'h21773321155;
assign testcases[7] = 44'h41851310064;
assign testcases[8] = 44'h32881221055;
assign testcases[9] = 44'h55895426644;
assign testcases[10] = 44'h22773321153;
assign testcases[11] = 44'h55895426644;
assign testcases[12] = 44'h42b53321051;
assign testcases[13] = 44'h2c791231555;
assign testcases[14] = 44'h255a8b43356;
assign testcases[15] = 44'h265a8b43356;
assign testcases[16] = 44'h54785821926;
assign testcases[17] = 44'h295833a1455;
assign testcases[18] = 44'h12891124154;
assign testcases[19] = 44'h27483491825;
assign testcases[20] = 44'h22883621816;
assign testcases[21] = 44'h33aa4522534;
assign testcases[22] = 44'h36582231335;
assign testcases[23] = 44'h22583222246;
assign testcases[24] = 44'h33982522233;
assign testcases[25] = 44'h22861221332;
assign testcases[26] = 44'h32770121434;
assign testcases[27] = 44'h36582231335;
assign testcases[28] = 44'h22982321064;
assign testcases[29] = 44'h32871221065;
assign testcases[30] = 44'h42874422163;
assign testcases[31] = 44'h52982522063;
assign testcases[32] = 44'h33586322265;
assign testcases[33] = 44'h229b492b253;
assign testcases[34] = 44'h22872321421;
assign testcases[35] = 44'h328a1125065;
assign testcases[36] = 44'h63991022255;
assign testcases[37] = 44'h34681311435;
assign testcases[38] = 44'h31a511411b2;
assign testcases[39] = 44'h55795225644;
assign testcases[40] = 44'h55795225644;
assign testcases[41] = 44'h22792422556;
assign testcases[42] = 44'h55680292344;
assign testcases[43] = 44'h58781221465;
assign testcases[44] = 44'h32970111063;
assign testcases[45] = 44'hc2f43211240;
assign testcases[46] = 44'h24686531794;
assign testcases[47] = 44'h32682231826;
assign testcases[48] = 44'h22870111433;
assign testcases[49] = 44'h22765221621;
assign testcases[50] = 44'h24581121466;
assign testcases[51] = 44'h23861221143;
assign testcases[52] = 44'h23860111143;
assign testcases[53] = 44'h22686722636;
assign testcases[54] = 44'h43564732244;
assign testcases[55] = 44'h32892523154;
assign testcases[56] = 44'h33480123938;
assign testcases[57] = 44'h247a6b35264;
assign testcases[58] = 44'h42993422355;
assign testcases[59] = 44'h22872222534;
assign testcases[60] = 44'h23993421636;
assign testcases[61] = 44'h24686431864;
assign testcases[62] = 44'h33882221344;
assign testcases[63] = 44'h32883321173;
assign testcases[64] = 44'h61870124174;
assign testcases[65] = 44'h61870124174;
assign testcases[66] = 44'h32982221244;
assign testcases[67] = 44'h62971121163;
assign testcases[68] = 44'h64783621927;
assign testcases[69] = 44'h56871221165;
assign testcases[70] = 44'h32781321164;
assign testcases[71] = 44'h31775421464;
assign testcases[72] = 44'h31775421464;
assign testcases[73] = 44'h22792221465;
assign testcases[74] = 44'h357a4622927;
assign testcases[75] = 44'h53aa2221a36;
assign testcases[76] = 44'h53aa2221a36;
assign testcases[77] = 44'h62a81322073;
assign testcases[78] = 44'h42874221273;
assign testcases[79] = 44'h28586621365;
assign testcases[80] = 44'h22871021342;
assign testcases[81] = 44'h295935c1b35;
assign testcases[82] = 44'h22884521844;
assign testcases[83] = 44'h285833a1464;
assign testcases[84] = 44'h54973421822;
assign testcases[85] = 44'h42872421253;
assign testcases[86] = 44'h4f287431446;
assign testcases[87] = 44'h33881211444;
assign testcases[88] = 44'h39597731737;
assign testcases[89] = 44'h12991221153;
assign testcases[90] = 44'h32678921445;
assign testcases[91] = 44'h4f287431446;
assign testcases[92] = 44'h3f287431546;
assign testcases[93] = 44'h33881211444;
assign testcases[94] = 44'h51d449111a1;
assign testcases[95] = 44'hb3e46412350;
assign testcases[96] = 44'h62981222073;
assign testcases[97] = 44'h23671021443;
assign testcases[98] = 44'h32880122194;
assign testcases[99] = 44'h12782321355;
assign testcases[100] = 44'h43882221555;
assign testcases[101] = 44'h52771221545;
assign testcases[102] = 44'h12782321355;
assign testcases[103] = 44'h22783221455;
assign testcases[104] = 44'h21772121444;
assign testcases[105] = 44'h22783221455;
assign testcases[106] = 44'h294844c1b35;
assign testcases[107] = 44'h24983321562;
assign testcases[108] = 44'h35894422825;
assign testcases[109] = 44'h23688831875;
assign testcases[110] = 44'h36672221355;
assign testcases[111] = 44'h33576221155;
assign testcases[112] = 44'h33576321255;
assign testcases[113] = 44'h337a2522728;
assign testcases[114] = 44'h36672221355;
assign testcases[115] = 44'h53483321537;
assign testcases[116] = 44'h43892221455;
assign testcases[117] = 44'h22881121255;
assign testcases[118] = 44'h63673331156;
assign testcases[119] = 44'h22875521163;
assign testcases[120] = 44'h127752411a4;
assign testcases[121] = 44'h63673331156;
assign testcases[122] = 44'h22990022064;
assign testcases[123] = 44'h32992222065;
assign testcases[124] = 44'h31875521345;
assign testcases[125] = 44'h245a5641156;
assign testcases[126] = 44'h62a700210d5;
assign testcases[127] = 44'h61a700210d5;
assign testcases[128] = 44'h56971011355;
assign testcases[129] = 44'h22961121232;
assign testcases[130] = 44'h23687731975;
assign testcases[131] = 44'hb3b45412141;
assign testcases[132] = 44'hb3b45412141;
assign testcases[133] = 44'h32861411043;
assign testcases[134] = 44'h426713211a5;
assign testcases[135] = 44'h35683321275;
assign testcases[136] = 44'h34683221275;
assign testcases[137] = 44'h23982321634;
assign testcases[138] = 44'h32776321355;
assign testcases[139] = 44'h32776421355;
assign testcases[140] = 44'h35683321275;
assign testcases[141] = 44'h34683221275;
assign testcases[142] = 44'he4c23611021;
assign testcases[143] = 44'h22861011132;
assign testcases[144] = 44'he4c23611021;
assign testcases[145] = 44'h23588731965;
assign testcases[146] = 44'h42a55521062;
assign testcases[147] = 44'h25585261444;
assign testcases[148] = 44'h42971222243;
assign testcases[149] = 44'h53a92222735;
assign testcases[150] = 44'h52770121824;
assign testcases[151] = 44'h2f0b47f3f47;
assign testcases[152] = 44'h42865521054;
assign testcases[153] = 44'h42865521054;
assign testcases[154] = 44'h54987625734;
assign testcases[155] = 44'h54987625734;
assign testcases[156] = 44'h54987625734;
assign testcases[157] = 44'h54987625734;
assign testcases[158] = 44'h22981221064;
assign testcases[159] = 44'h22b85421353;
assign testcases[160] = 44'h32671121094;
assign testcases[161] = 44'h27581220064;
assign testcases[162] = 44'h42771421145;
assign testcases[163] = 44'h228a7827454;
assign testcases[164] = 44'h22897827454;
assign testcases[165] = 44'h33675321865;
assign testcases[166] = 44'h42865421263;
assign testcases[167] = 44'h11862421054;
assign testcases[168] = 44'h52962221163;
assign testcases[169] = 44'h3c373391464;
assign testcases[170] = 44'h20880111085;
assign testcases[171] = 44'h23781121335;
assign testcases[172] = 44'h23781121335;
assign testcases[173] = 44'h82972511154;
assign testcases[174] = 44'h31772121334;
assign testcases[175] = 44'h34872421143;
assign testcases[176] = 44'h31772121334;
assign testcases[177] = 44'h53b82222744;
assign testcases[178] = 44'h32981112083;
assign testcases[179] = 44'h32682212256;
assign testcases[180] = 44'h32682212256;
assign testcases[181] = 44'h27586571856;
assign testcases[182] = 44'h22982322074;
assign testcases[183] = 44'h22a83221353;
assign testcases[184] = 44'h22a83221353;
assign testcases[185] = 44'h32784631926;
assign testcases[186] = 44'h22883321834;
assign testcases[187] = 44'h32891222264;
assign testcases[188] = 44'h32688321545;
assign testcases[189] = 44'h32688421545;
assign testcases[190] = 44'h23697522645;
assign testcases[191] = 44'h33a92521433;
assign testcases[192] = 44'h33787323263;
assign testcases[193] = 44'h32771121354;
assign testcases[194] = 44'h32771121354;
assign testcases[195] = 44'h22686521555;
assign testcases[196] = 44'h42983322554;
assign testcases[197] = 44'h46591211a2a;
assign testcases[198] = 44'hb5a35310181;
assign testcases[199] = 44'h71a612111b3;
assign testcases[200] = 44'h55681211827;
assign testcases[201] = 44'h27498921836;
assign testcases[202] = 44'h34862321243;
assign testcases[203] = 44'h22872321633;
assign testcases[204] = 44'h22872321633;
assign testcases[205] = 44'h646b1222c2c;
assign testcases[206] = 44'h646b1222c2c;
assign testcases[207] = 44'h22776621555;
assign testcases[208] = 44'h23685422445;
assign testcases[209] = 44'h55791111929;
assign testcases[210] = 44'ha5771111a47;
assign testcases[211] = 44'h42883222475;
assign testcases[212] = 44'h43691111a4a;
assign testcases[213] = 44'h41773611455;
assign testcases[214] = 44'h34692222175;
assign testcases[215] = 44'h54897615843;
assign testcases[216] = 44'h62572321366;
assign testcases[217] = 44'h22882221475;
assign testcases[218] = 44'h32872221344;
assign testcases[219] = 44'h33788522545;
assign testcases[220] = 44'h22873521625;
assign testcases[221] = 44'h22574321444;
assign testcases[222] = 44'h33960111153;
assign testcases[223] = 44'h43791221466;
assign testcases[224] = 44'h52793321665;
assign testcases[225] = 44'h52873622434;
assign testcases[226] = 44'h3c474691856;
assign testcases[227] = 44'h338a1222286;
assign testcases[228] = 44'h52873622434;
assign testcases[229] = 44'h62982222443;
assign testcases[230] = 44'h93a36411141;
assign testcases[231] = 44'h42872221135;
assign testcases[232] = 44'h34893422336;
assign testcases[233] = 44'h62982222443;
assign testcases[234] = 44'h127821121a5;
assign testcases[235] = 44'h12882321064;
assign testcases[236] = 44'h12882321064;
assign testcases[237] = 44'h22882321064;
assign testcases[238] = 44'h12882321064;
assign testcases[239] = 44'h127821121a5;
assign testcases[240] = 44'h27383171666;
assign testcases[241] = 44'h645b112193a;
assign testcases[242] = 44'h32476621254;
assign testcases[243] = 44'h254c122171f;
assign testcases[244] = 44'h254c122171f;
assign testcases[245] = 44'h46ba1121064;
assign testcases[246] = 44'h32883321164;
assign testcases[247] = 44'h21674222355;
assign testcases[248] = 44'h31872221144;
assign testcases[249] = 44'h46ba1121064;
assign testcases[250] = 44'h446a2311729;
assign testcases[251] = 44'h44982321054;
assign testcases[252] = 44'h525a1122839;
assign testcases[253] = 44'h32675221774;
assign testcases[254] = 44'h44982321054;
assign testcases[255] = 44'h22786423455;
assign testcases[256] = 44'h23690121627;
assign testcases[257] = 44'h23983221063;
assign testcases[258] = 44'h294822f1c34;
assign testcases[259] = 44'h558b2322828;
assign testcases[260] = 44'h23772421425;
assign testcases[261] = 44'h23873221193;
assign testcases[262] = 44'h42872221045;
assign testcases[263] = 44'h23772521435;
assign testcases[264] = 44'h654c111285b;
assign testcases[265] = 44'h4468012182a;
assign testcases[266] = 44'h34bc3623085;
assign testcases[267] = 44'hb5882323735;
assign testcases[268] = 44'h26ca1122153;
assign testcases[269] = 44'h467b112381a;
assign testcases[270] = 44'h63883623155;
assign testcases[271] = 44'h467b112381a;
assign testcases[272] = 44'h446b3423939;
assign testcases[273] = 44'h23792222375;
assign testcases[274] = 44'h248b5627364;
assign testcases[275] = 44'h63883623155;
assign testcases[276] = 44'h26ca1122153;
assign testcases[277] = 44'h467b112381a;
assign testcases[278] = 44'ha5690126728;
assign testcases[279] = 44'h548b2225536;
assign testcases[280] = 44'h255a112372a;
assign testcases[281] = 44'h47680193b24;
assign testcases[282] = 44'h22883212244;
assign testcases[283] = 44'h548b2225536;
assign testcases[284] = 44'h347c4723158;
assign testcases[285] = 44'h347c4723158;
assign testcases[286] = 44'h545b252194a;
assign testcases[287] = 44'h54883622234;
assign testcases[288] = 44'h55892422146;
assign testcases[289] = 44'h266d572383a;
assign testcases[290] = 44'h55892422146;
assign testcases[291] = 44'h54791191819;
assign testcases[292] = 44'h536b2422458;
assign testcases[293] = 44'h43871122433;
assign testcases[294] = 44'h354d342382c;
assign testcases[295] = 44'h334c1122749;
assign testcases[296] = 44'h42594622688;
assign testcases[297] = 44'h34ca1221164;
assign testcases[298] = 44'h35cb1122064;
assign testcases[299] = 44'h34ca2221163;
assign testcases[300] = 44'h62882422144;
assign testcases[301] = 44'h43681111819;
assign testcases[302] = 44'h44ab1222265;
assign testcases[303] = 44'h32871151264;
assign testcases[304] = 44'h22685231a65;
assign testcases[305] = 44'h225b1112848;
assign testcases[306] = 44'h22883121554;
assign testcases[307] = 44'h336b0152738;
assign testcases[308] = 44'h336b0152738;
assign testcases[309] = 44'h32881211624;
assign testcases[310] = 44'h225b1112848;
assign testcases[311] = 44'h22776321445;
assign testcases[312] = 44'h33795422546;
assign testcases[313] = 44'h22797722546;
assign testcases[314] = 44'h63874622534;
assign testcases[315] = 44'h63973422534;
assign testcases[316] = 44'h437b5823457;
assign testcases[317] = 44'h537a4722277;
assign testcases[318] = 44'h848a3523667;
assign testcases[319] = 44'h537a4722277;
assign testcases[320] = 44'h848a3523667;
assign testcases[321] = 44'h336b5523457;
assign testcases[322] = 44'h23791122155;
assign testcases[323] = 44'h347a4822758;
assign testcases[324] = 44'h235d232b348;
assign testcases[325] = 44'h235d232b348;
assign testcases[326] = 44'h84490133b4a;
assign testcases[327] = 44'h85790134848;
assign testcases[328] = 44'h335c1122a2c;
assign testcases[329] = 44'h33691111649;
assign testcases[330] = 44'ha3692232a38;
assign testcases[331] = 44'ha3692232a38;
assign testcases[332] = 44'h22686513455;
assign testcases[333] = 44'h62572321155;
assign testcases[334] = 44'h84872422065;
assign testcases[335] = 44'h955b113386a;
assign testcases[336] = 44'ha4861111736;
assign testcases[337] = 44'h53793622535;
assign testcases[338] = 44'h865d562294b;
assign testcases[339] = 44'h3a5b122292b;
assign testcases[340] = 44'h285c121282b;
assign testcases[341] = 44'h75681112838;
assign testcases[342] = 44'h347a0131839;
assign testcases[343] = 44'h347a0131839;
assign testcases[344] = 44'h645c112285a;
assign testcases[345] = 44'h45b93911063;
assign testcases[346] = 44'ha5b62422083;
assign testcases[347] = 44'h964a1122b4d;
assign testcases[348] = 44'h46592322557;
assign testcases[349] = 44'h258b1222076;
assign testcases[350] = 44'h467c2432469;
assign testcases[351] = 44'h258b1222076;
assign testcases[352] = 44'h24791222064;
assign testcases[353] = 44'hb46e4534d4d;
assign testcases[354] = 44'h92619911612;
assign testcases[355] = 44'hb3a61422073;
assign testcases[356] = 44'h657c362283a;
assign testcases[357] = 44'h84681232b38;
assign testcases[358] = 44'h555c1232b3a;
assign testcases[359] = 44'h335d2222b3b;
assign testcases[360] = 44'h24684321465;
assign testcases[361] = 44'h468a2522546;
assign testcases[362] = 44'h424b2122b5a;
assign testcases[363] = 44'h453a1121a4b;
assign testcases[364] = 44'h444e2125b5c;
assign testcases[365] = 44'h86791133838;
assign testcases[366] = 44'h444e2125b5c;
assign testcases[367] = 44'h135c1222a58;
assign testcases[368] = 44'h236b4342828;
assign testcases[369] = 44'h98671122827;
assign testcases[370] = 44'h44a93812073;
assign testcases[371] = 44'h15781211615;
assign testcases[372] = 44'h57782611826;
assign testcases[373] = 44'h23474231454;
assign testcases[374] = 44'h653d2123a3d;
assign testcases[375] = 44'h853a1134b5a;
assign testcases[376] = 44'h677c242284a;
assign testcases[377] = 44'h98671122827;
assign testcases[378] = 44'hc65a1126b6a;
assign testcases[379] = 44'h64793522635;
assign testcases[380] = 44'h25691221725;
assign testcases[381] = 44'h454d2422b3d;
assign testcases[382] = 44'h25691221725;
assign testcases[383] = 44'h25691221725;
assign testcases[384] = 44'h24993521444;
assign testcases[385] = 44'h34992222164;
assign testcases[386] = 44'h24892521455;
assign testcases[387] = 44'h32782421265;
assign testcases[388] = 44'h24993521445;
assign testcases[389] = 44'h446a2322537;
assign testcases[390] = 44'hb5a35211181;
assign testcases[391] = 44'h454d2422b3d;
assign testcases[392] = 44'h32691121837;
assign testcases[393] = 44'h22585331a65;
assign testcases[394] = 44'h424b1112a5b;
assign testcases[395] = 44'hb36c2114c3a;
assign testcases[396] = 44'h429b7f38073;
assign testcases[397] = 44'h636a232295a;
assign testcases[398] = 44'h636a232295a;
assign testcases[399] = 44'h22572212476;
assign testcases[400] = 44'h429b7f38073;
assign testcases[401] = 44'h61762411524;
assign testcases[402] = 44'h535c342294b;
assign testcases[403] = 44'h535b222285a;
assign testcases[404] = 44'h23791322164;
assign testcases[405] = 44'h44881211726;
assign testcases[406] = 44'h63691212847;
assign testcases[407] = 44'h636b1222b3a;
assign testcases[408] = 44'h74681143928;
assign testcases[409] = 44'h3249262484b;
assign testcases[410] = 44'h338a5622536;
assign testcases[411] = 44'h338a4522646;
assign testcases[412] = 44'h23784321374;
assign testcases[413] = 44'h857a1126838;
assign testcases[414] = 44'h337a7522546;
assign testcases[415] = 44'h277d7736476;
assign testcases[416] = 44'h83781131a48;
assign testcases[417] = 44'h51967721253;
assign testcases[418] = 44'h546b113183a;
assign testcases[419] = 44'h43b93711073;
assign testcases[420] = 44'h84783822557;
assign testcases[421] = 44'ha2a62712083;
assign testcases[422] = 44'h61863311394;
assign testcases[423] = 44'h65591111818;
assign testcases[424] = 44'h61863311394;
assign testcases[425] = 44'ha2a62712083;
assign testcases[426] = 44'h72962411163;
assign testcases[427] = 44'h527a1121477;
assign testcases[428] = 44'h23691220546;
assign testcases[429] = 44'h535b2322a8c;
assign testcases[430] = 44'h65591111818;
assign testcases[431] = 44'h22693521655;
assign testcases[432] = 44'hb3371222b3a;
assign testcases[433] = 44'h325c1122a3b;
assign testcases[434] = 44'h455b3523938;
assign testcases[435] = 44'h325c1122a3b;
assign testcases[436] = 44'h42773811565;
assign testcases[437] = 44'h735a1113c49;
assign testcases[438] = 44'h455b3523938;
assign testcases[439] = 44'h23462111353;
assign testcases[440] = 44'h352a1121c2b;
assign testcases[441] = 44'h734a1111a3a;
assign testcases[442] = 44'h733f2123c6f;
assign testcases[443] = 44'h83671222848;
assign testcases[444] = 44'ha5a41111051;
assign testcases[445] = 44'h426a1121277;
assign testcases[446] = 44'h545b4722a3b;
assign testcases[447] = 44'h74681131547;
assign testcases[448] = 44'h42681121446;
assign testcases[449] = 44'h635b2422b3a;
assign testcases[450] = 44'h635b2422b3a;
assign testcases[451] = 44'h274912b1835;
assign testcases[452] = 44'h43982421053;
assign testcases[453] = 44'h747b1122a28;
assign testcases[454] = 44'h73a63511613;
assign testcases[455] = 44'hc36a1125b59;
assign testcases[456] = 44'h528a1122656;
assign testcases[457] = 44'h327a3622367;
assign testcases[458] = 44'h747b1122a28;
assign testcases[459] = 44'h126d2221b5a;
assign testcases[460] = 44'h73891322837;
assign testcases[461] = 44'h237a1122455;
assign testcases[462] = 44'h83681222b29;
assign testcases[463] = 44'h12487521b65;
assign testcases[464] = 44'h243a112192a;
assign testcases[465] = 44'h369c1222628;
assign testcases[466] = 44'h845a3521748;
assign testcases[467] = 44'he4751112746;
assign testcases[468] = 44'h235c1121b3a;
assign testcases[469] = 44'h32662820086;
assign testcases[470] = 44'h534b2322a2c;
assign testcases[471] = 44'h74683522757;
assign testcases[472] = 44'h555b452293b;
assign testcases[473] = 44'h54780111938;
assign testcases[474] = 44'h256a1221828;
assign testcases[475] = 44'h435a1121467;
assign testcases[476] = 44'h34791121727;
assign testcases[477] = 44'h67691121818;
assign testcases[478] = 44'h435a1121467;
assign testcases[479] = 44'h446a1122267;
assign testcases[480] = 44'h235f112f628;
assign testcases[481] = 44'h86571122927;
assign testcases[482] = 44'h274a1141938;
assign testcases[483] = 44'h274a1141a38;
assign testcases[484] = 44'hc3481134b48;
assign testcases[485] = 44'h41591111668;
assign testcases[486] = 44'h41591111668;
assign testcases[487] = 44'h415a0111668;
assign testcases[488] = 44'h667c382292a;
assign testcases[489] = 44'h448a1222637;
assign testcases[490] = 44'h537a3522477;
assign testcases[491] = 44'hc4861212837;
assign testcases[492] = 44'hc5761312836;
assign testcases[493] = 44'h849c4522566;
assign testcases[494] = 44'h92965618433;
assign testcases[495] = 44'h63581122839;
assign testcases[496] = 44'h139a2321445;
assign testcases[497] = 44'h74786922524;
assign testcases[498] = 44'h63581122839;
assign testcases[499] = 44'h849c4522566;
assign testcases[500] = 44'h139a2321445;
assign testcases[501] = 44'h955a4826c48;
assign testcases[502] = 44'h955a4826c48;
assign testcases[503] = 44'h67691121828;
assign testcases[504] = 44'h67691121718;
assign testcases[505] = 44'ha4581222a48;
assign testcases[506] = 44'h67691121718;
assign testcases[507] = 44'h345c0122969;
assign testcases[508] = 44'h436b3621558;
assign testcases[509] = 44'h734a2522c2c;
assign testcases[510] = 44'h3349242483b;
assign testcases[511] = 44'h436b3621558;
assign testcases[512] = 44'h35492331839;
assign testcases[513] = 44'h83481132a48;
assign testcases[514] = 44'h83481132a48;
assign testcases[515] = 44'h287d8736866;
assign testcases[516] = 44'h946d012485b;
assign testcases[517] = 44'h035b1151858;
assign testcases[518] = 44'h83681222819;
assign testcases[519] = 44'h64886922834;
assign testcases[520] = 44'h459a2322817;
assign testcases[521] = 44'h23992321834;
assign testcases[522] = 44'h36897a22835;
assign testcases[523] = 44'h22698822837;
assign testcases[524] = 44'h33696522837;
assign testcases[525] = 44'h436b3622468;
assign testcases[526] = 44'h64886922834;
assign testcases[527] = 44'h74874722833;
assign testcases[528] = 44'h148a3722835;
assign testcases[529] = 44'h22492122468;
assign testcases[530] = 44'h558a1021416;
assign testcases[531] = 44'h535c222283a;
assign testcases[532] = 44'h535c222283a;
assign testcases[533] = 44'hb3662321428;
assign testcases[534] = 44'h427c1322448;
assign testcases[535] = 44'h558a1021416;
assign testcases[536] = 44'h22492122468;
assign testcases[537] = 44'h64880121485;
assign testcases[538] = 44'h936d211583c;
assign testcases[539] = 44'h736b1125c49;
assign testcases[540] = 44'h337a2423457;
assign testcases[541] = 44'h646a1116847;
assign testcases[542] = 44'h42581121477;
assign testcases[543] = 44'h644b3322469;
assign testcases[544] = 44'h042d1121c2e;
assign testcases[545] = 44'h224a6822846;
assign testcases[546] = 44'h349a1221454;
assign testcases[547] = 44'h657a1112828;
assign testcases[548] = 44'h545b462283b;
assign testcases[549] = 44'h23791141846;
assign testcases[550] = 44'h32771221043;
assign testcases[551] = 44'h44692322437;
assign testcases[552] = 44'h44592322447;
assign testcases[553] = 44'h83d457114a1;
assign testcases[554] = 44'h742f122486f;
assign testcases[555] = 44'h742f122486f;
assign testcases[556] = 44'h824c1234849;
assign testcases[557] = 44'h742f122486f;
assign testcases[558] = 44'h824c1234849;
assign testcases[559] = 44'hb37e212484c;
assign testcases[560] = 44'h725b112285b;
assign testcases[561] = 44'h22697622846;
assign testcases[562] = 44'h234a6922856;
assign testcases[563] = 44'h43783522824;
assign testcases[564] = 44'hb37e212484c;
assign testcases[565] = 44'h725b112285b;
assign testcases[566] = 44'h137b1162466;
assign testcases[567] = 44'h137b1162466;
assign testcases[568] = 44'h647a1162847;
assign testcases[569] = 44'h82a52421432;
assign testcases[570] = 44'h667c222383a;
assign testcases[571] = 44'h82a52421432;
assign testcases[572] = 44'h53591222818;
assign testcases[573] = 44'h327b2321858;
assign testcases[574] = 44'h446b4423828;
assign testcases[575] = 44'h456b262282b;
assign testcases[576] = 44'h42890122448;
assign testcases[577] = 44'h337a6422846;
assign testcases[578] = 44'h337a6422846;
assign testcases[579] = 44'h32592411828;
assign testcases[580] = 44'h316c012184b;
assign testcases[581] = 44'h316c012184b;
assign testcases[582] = 44'h216c112184a;
assign testcases[583] = 44'h4339122182a;
assign testcases[584] = 44'h647c4c2382a;
assign testcases[585] = 44'h33992222444;
assign testcases[586] = 44'h575a2322829;
assign testcases[587] = 44'h22785431474;
assign testcases[588] = 44'he4c22411431;
assign testcases[589] = 44'h54490112828;
assign testcases[590] = 44'h328a4522846;
assign testcases[591] = 44'h82538521833;
assign testcases[592] = 44'h328a4522846;
assign testcases[593] = 44'h127c2223948;
assign testcases[594] = 44'h32892422375;
assign testcases[595] = 44'h227b6728756;
assign testcases[596] = 44'h234b111183b;
assign testcases[597] = 44'h4349112195a;
assign testcases[598] = 44'h31681121356;
assign testcases[599] = 44'h243c122275b;
assign testcases[600] = 44'h41771121495;
assign testcases[601] = 44'h125c222184c;
assign testcases[602] = 44'h22790122084;
assign testcases[603] = 44'h125c222184c;
assign testcases[604] = 44'h235a3322255;
assign testcases[605] = 44'h227a1122255;
assign testcases[606] = 44'h94881224837;
assign testcases[607] = 44'h527a3623746;
assign testcases[608] = 44'h537f3235668;
assign testcases[609] = 44'hb2a62323332;
assign testcases[610] = 44'h228a3522916;
assign testcases[611] = 44'h223c112293c;
assign testcases[612] = 44'h43781422064;
assign testcases[613] = 44'h34771211635;
assign testcases[614] = 44'h4a285241377;
assign testcases[615] = 44'h32ab4622857;
assign testcases[616] = 44'h32ab4622857;
assign testcases[617] = 44'h364a132182a;
assign testcases[618] = 44'h445c113284a;
assign testcases[619] = 44'h254a1122739;
assign testcases[620] = 44'h23796323455;
assign testcases[621] = 44'h23796323455;
assign testcases[622] = 44'h32591221458;
assign testcases[623] = 44'h96992522445;
assign testcases[624] = 44'h449b3535063;
assign testcases[625] = 44'h449b3535063;
assign testcases[626] = 44'h228a1121556;
assign testcases[627] = 44'h228a1121556;
assign testcases[628] = 44'h23791122456;
assign testcases[629] = 44'h23674432464;
assign testcases[630] = 44'h23791122456;
assign testcases[631] = 44'h336a1122928;
assign testcases[632] = 44'h52772522234;
assign testcases[633] = 44'h739d5223498;
assign testcases[634] = 44'h32775a21335;
assign testcases[635] = 44'h32762511086;
assign testcases[636] = 44'h22698722487;
assign testcases[637] = 44'h22698722487;
assign testcases[638] = 44'h43871131294;
assign testcases[639] = 44'h5a683511626;
assign testcases[640] = 44'h238b2322758;
assign testcases[641] = 44'h339b4522757;
assign testcases[642] = 44'h238b2322758;
assign testcases[643] = 44'h339b4522757;
assign testcases[644] = 44'h238b2322758;
assign testcases[645] = 44'h438a0136265;
assign testcases[646] = 44'h43881133164;
assign testcases[647] = 44'h62780121085;
assign testcases[648] = 44'h73771212546;
assign testcases[649] = 44'h72568518433;
assign testcases[650] = 44'h322a1231639;
assign testcases[651] = 44'h738d8822487;
assign testcases[652] = 44'hf5394527a3f;
assign testcases[653] = 44'h92591222927;
assign testcases[654] = 44'h31491122846;
assign testcases[655] = 44'h235c3422357;
assign testcases[656] = 44'h322a1231639;
assign testcases[657] = 44'h5329252194a;
assign testcases[658] = 44'h35781121144;
assign testcases[659] = 44'h62880124084;
assign testcases[660] = 44'h35781121144;
assign testcases[661] = 44'h13792321534;
assign testcases[662] = 44'h34881221154;
assign testcases[663] = 44'h44490111728;
assign testcases[664] = 44'h434c332183b;
assign testcases[665] = 44'h32592521257;
assign testcases[666] = 44'h33691161645;
assign testcases[667] = 44'h233a1121729;
assign testcases[668] = 44'h62581312778;
assign testcases[669] = 44'h233a1121729;
assign testcases[670] = 44'h42772722433;
assign testcases[671] = 44'h32680121375;
assign testcases[672] = 44'h325987215c7;
assign testcases[673] = 44'h32680121375;
assign testcases[674] = 44'h234a1121739;
assign testcases[675] = 44'h437a1211637;
assign testcases[676] = 44'h234a1121739;
assign testcases[677] = 44'h41891222276;
assign testcases[678] = 44'h429a5a22275;
assign testcases[679] = 44'h32582413729;
assign testcases[680] = 44'h124c232193c;
assign testcases[681] = 44'h42671321445;
assign testcases[682] = 44'h32793721546;
assign testcases[683] = 44'h72881112475;
assign testcases[684] = 44'h21698822597;
assign testcases[685] = 44'h72881112475;
assign testcases[686] = 44'h23982321364;
assign testcases[687] = 44'h327b2322466;
assign testcases[688] = 44'h21870111164;
assign testcases[689] = 44'h27791141835;
assign testcases[690] = 44'h62b801240c4;
assign testcases[691] = 44'h329b5222497;
assign testcases[692] = 44'h184933b1846;
assign testcases[693] = 44'h237a7522546;
assign testcases[694] = 44'h237a7522546;
assign testcases[695] = 44'hb3f22410041;
assign testcases[696] = 44'h33981211063;
assign testcases[697] = 44'h33981211063;
assign testcases[698] = 44'h327c4423457;
assign testcases[699] = 44'h635a112193a;
assign testcases[700] = 44'h424a56227a8;
assign testcases[701] = 44'h33981211063;
assign testcases[702] = 44'h23981211063;
assign testcases[703] = 44'h34784522834;
assign testcases[704] = 44'h32790121176;
assign testcases[705] = 44'h428a32262a5;
assign testcases[706] = 44'h41861221173;
assign testcases[707] = 44'h52882322344;
assign testcases[708] = 44'h83872212255;
assign testcases[709] = 44'h437a2311827;
assign testcases[710] = 44'h424a45227a8;
assign testcases[711] = 44'h338b6322556;
assign testcases[712] = 44'h218b2323066;
assign testcases[713] = 44'h21892222635;
assign testcases[714] = 44'h32794522478;
assign testcases[715] = 44'h21782322344;
assign testcases[716] = 44'h21892222635;
assign testcases[717] = 44'h42682222244;
assign testcases[718] = 44'h31691221155;
assign testcases[719] = 44'h32992423064;
assign testcases[720] = 44'h31691221155;
assign testcases[721] = 44'h225a6822446;
assign testcases[722] = 44'h42682322134;
assign testcases[723] = 44'h3c387811524;
assign testcases[724] = 44'h73a701222b4;
assign testcases[725] = 44'h52790122366;
assign testcases[726] = 44'h749b2422175;
assign testcases[727] = 44'h33980111053;
assign testcases[728] = 44'h33980111053;
assign testcases[729] = 44'hb2b63623083;
assign testcases[730] = 44'h335a22a2b57;
assign testcases[731] = 44'h829b0123286;
assign testcases[732] = 44'h31881221084;
assign testcases[733] = 44'h33a94322543;
assign testcases[734] = 44'h239a2221354;
assign testcases[735] = 44'h32771231294;
assign testcases[736] = 44'h32771231294;
assign testcases[737] = 44'h23ac3422055;
assign testcases[738] = 44'h225a6622446;
assign testcases[739] = 44'h238a2422066;
assign testcases[740] = 44'h83981224575;
assign testcases[741] = 44'h32698622447;
assign testcases[742] = 44'h23981211053;
assign testcases[743] = 44'h425c552293a;
assign testcases[744] = 44'h325c5522939;
assign testcases[745] = 44'h34a91221344;
assign testcases[746] = 44'h11793222625;
assign testcases[747] = 44'h21794322626;
assign testcases[748] = 44'h34a91221344;
assign testcases[749] = 44'h34a91221344;
assign testcases[750] = 44'h32792422265;
assign testcases[751] = 44'h32792422265;
assign testcases[752] = 44'h23893522254;
assign testcases[753] = 44'h32792422265;
assign testcases[754] = 44'h274813b1b45;
assign testcases[755] = 44'h61a62511195;
assign testcases[756] = 44'h71b62311092;
assign testcases[757] = 44'h32681221085;
assign testcases[758] = 44'h32681221085;
assign testcases[759] = 44'h226a5722336;
assign testcases[760] = 44'h32696222456;
assign testcases[761] = 44'h31692121467;
assign testcases[762] = 44'h42781221066;
assign testcases[763] = 44'h31692121467;
assign testcases[764] = 44'h327a2222266;
assign testcases[765] = 44'h327a2222267;
assign testcases[766] = 44'h22594222356;
assign testcases[767] = 44'h339b5322554;
assign testcases[768] = 44'h32a95522054;
assign testcases[769] = 44'h32881121075;
assign testcases[770] = 44'h32a95522054;
assign testcases[771] = 44'h22798522467;
assign testcases[772] = 44'h22798522457;
assign testcases[773] = 44'h36782041535;
assign testcases[774] = 44'h36782041535;
assign testcases[775] = 44'h419711220a4;
assign testcases[776] = 44'h53872162373;
assign testcases[777] = 44'h52871162363;
assign testcases[778] = 44'h53892123535;
assign testcases[779] = 44'h33a95522044;
assign testcases[780] = 44'h23782251053;
assign testcases[781] = 44'h33c92232243;
assign testcases[782] = 44'h42895622186;
assign testcases[783] = 44'h33c92232243;
assign testcases[784] = 44'h32a94422054;
assign testcases[785] = 44'h326a3222738;
assign testcases[786] = 44'h326a3222738;
assign testcases[787] = 44'h426b3421458;
assign testcases[788] = 44'h426b3421458;
assign testcases[789] = 44'h22496522366;
assign testcases[790] = 44'h33784422734;
assign testcases[791] = 44'h326a7522366;
assign testcases[792] = 44'h33995422054;
assign testcases[793] = 44'h62870112054;
assign testcases[794] = 44'ha2561112928;
assign testcases[795] = 44'h48393132589;
assign testcases[796] = 44'h34593532546;
assign testcases[797] = 44'h65662511737;
assign testcases[798] = 44'h627a0123547;
assign testcases[799] = 44'h627a0123547;
assign testcases[800] = 44'h22676623154;
assign testcases[801] = 44'h41691213156;
assign testcases[802] = 44'hb6a35311051;
assign testcases[803] = 44'h33682332154;
assign testcases[804] = 44'h42781122445;
assign testcases[805] = 44'hb4740112625;
assign testcases[806] = 44'ha4740111615;
assign testcases[807] = 44'hb4740112625;
assign testcases[808] = 44'h25780141244;
assign testcases[809] = 44'h52681122544;
assign testcases[810] = 44'h51770112244;
assign testcases[811] = 44'h634c112294c;
assign testcases[812] = 44'h646a2422549;
assign testcases[813] = 44'h72950121433;
assign testcases[814] = 44'h746b242293b;
assign testcases[815] = 44'h646a2422549;
assign testcases[816] = 44'h526a1223347;
assign testcases[817] = 44'h94761421729;
assign testcases[818] = 44'h21772522074;
assign testcases[819] = 44'h327b3223266;
assign testcases[820] = 44'h33871221063;
assign testcases[821] = 44'he4c22311030;
assign testcases[822] = 44'h33b82321253;
assign testcases[823] = 44'h33b82321253;
assign testcases[824] = 44'h52681112444;
assign testcases[825] = 44'h62872322244;
assign testcases[826] = 44'h63860112524;
assign testcases[827] = 44'h62872322244;
assign testcases[828] = 44'hb4952712155;
assign testcases[829] = 44'h74a41321152;
assign testcases[830] = 44'h62870112164;
assign testcases[831] = 44'h74a41321152;
assign testcases[832] = 44'h458a2741748;
assign testcases[833] = 44'h458a384174a;
assign testcases[834] = 44'h21781321466;
assign testcases[835] = 44'h22883611264;
assign testcases[836] = 44'h81715802423;
assign testcases[837] = 44'h81715802423;
assign testcases[838] = 44'h75681221628;
assign testcases[839] = 44'h41981321142;
assign testcases[840] = 44'h94692222839;
assign testcases[841] = 44'h53971532063;
assign testcases[842] = 44'h64684732748;
assign testcases[843] = 44'h23775221664;
assign testcases[844] = 44'h55672611718;
assign testcases[845] = 44'h33b81321363;
assign testcases[846] = 44'h33b81321363;
assign testcases[847] = 44'h44a92221364;
assign testcases[848] = 44'h33b81321363;
assign testcases[849] = 44'h33b81221363;
assign testcases[850] = 44'h32781221737;
assign testcases[851] = 44'h32781221737;
assign testcases[852] = 44'h37697622535;
assign testcases[853] = 44'h64983921637;
assign testcases[854] = 44'h64983921637;
assign testcases[855] = 44'h84a60222074;
assign testcases[856] = 44'h64983921637;
assign testcases[857] = 44'h74872322525;
assign testcases[858] = 44'h5358141182a;
assign testcases[859] = 44'h75851321453;
assign testcases[860] = 44'h32a94322154;
assign testcases[861] = 44'h83c45311ba2;
assign testcases[862] = 44'h51671112534;
assign testcases[863] = 44'h32a94422154;
assign testcases[864] = 44'h32a94322154;
assign testcases[865] = 44'h32a95322164;
assign testcases[866] = 44'h75851322443;
assign testcases[867] = 44'h75851321443;
assign testcases[868] = 44'h75851321453;
assign testcases[869] = 44'h63972621064;
assign testcases[870] = 44'h82842711074;
assign testcases[871] = 44'h52a62821053;
assign testcases[872] = 44'h42972611434;
assign testcases[873] = 44'h72660111616;
assign testcases[874] = 44'h83580121738;
assign testcases[875] = 44'h84771132626;
assign testcases[876] = 44'h62860111044;
assign testcases[877] = 44'h82842711074;
assign testcases[878] = 44'h42694723356;
assign testcases[879] = 44'h32a95422154;
assign testcases[880] = 44'h42571221357;
assign testcases[881] = 44'h73962711074;
assign testcases[882] = 44'h94661352525;
assign testcases[883] = 44'h32a95422154;
assign testcases[884] = 44'h42694723356;
assign testcases[885] = 44'h538a1222276;
assign testcases[886] = 44'h537a1222276;
assign testcases[887] = 44'h94573612649;
assign testcases[888] = 44'h72963722053;
assign testcases[889] = 44'h236f5536599;
assign testcases[890] = 44'h42973721424;
assign testcases[891] = 44'h32a95322064;
assign testcases[892] = 44'h23691221448;
assign testcases[893] = 44'h32a95322064;
assign testcases[894] = 44'h32a95421064;
assign testcases[895] = 44'h62962622054;
assign testcases[896] = 44'ha4752422625;
assign testcases[897] = 44'h62962622054;
assign testcases[898] = 44'ha4752422625;
assign testcases[899] = 44'h629a01230a5;
assign testcases[900] = 44'h83872212626;
assign testcases[901] = 44'h63b92322264;
assign testcases[902] = 44'h63b92322264;
assign testcases[903] = 44'h62871216153;
assign testcases[904] = 44'h62871216153;
assign testcases[905] = 44'h32696322357;
assign testcases[906] = 44'h64874222454;
assign testcases[907] = 44'h82b60121052;
assign testcases[908] = 44'h62963722244;
assign testcases[909] = 44'h82740110624;
assign testcases[910] = 44'hc2670033837;
assign testcases[911] = 44'h636b0039726;
assign testcases[912] = 44'h93780112748;
assign testcases[913] = 44'h93770024737;
assign testcases[914] = 44'h82740110624;
assign testcases[915] = 44'h93760021626;
assign testcases[916] = 44'h63b53141371;
assign testcases[917] = 44'h438a2629533;
assign testcases[918] = 44'h64774721535;
assign testcases[919] = 44'h85862821255;
assign testcases[920] = 44'h52691222637;
assign testcases[921] = 44'h64774721535;
assign testcases[922] = 44'h85862821255;
assign testcases[923] = 44'h438a2629533;
assign testcases[924] = 44'h75661312446;
assign testcases[925] = 44'h65974c11616;
assign testcases[926] = 44'h45994b12517;
assign testcases[927] = 44'h22694221365;
assign testcases[928] = 44'h75661312446;
assign testcases[929] = 44'h94751213626;
assign testcases[930] = 44'h54c91221053;
assign testcases[931] = 44'h33992321054;
assign testcases[932] = 44'h32983621534;
assign testcases[933] = 44'h33992321054;
assign testcases[934] = 44'h54c91221053;
assign testcases[935] = 44'h84864412626;
assign testcases[936] = 44'h84864412626;
assign testcases[937] = 44'h5349112186a;
assign testcases[938] = 44'hb4842512634;
assign testcases[939] = 44'h72b50121342;
assign testcases[940] = 44'ha4861321827;
assign testcases[941] = 44'ha2661224828;
assign testcases[942] = 44'h436a3322638;
assign testcases[943] = 44'h336a2222547;
assign testcases[944] = 44'h93761223825;
assign testcases[945] = 44'h74571121748;
assign testcases[946] = 44'h96791224948;
assign testcases[947] = 44'ha3750121825;
assign testcases[948] = 44'h94861221706;
assign testcases[949] = 44'h94861221706;
assign testcases[950] = 44'h94861221706;
assign testcases[951] = 44'ha3750121825;
assign testcases[952] = 44'h73760111625;
assign testcases[953] = 44'h93650111828;
assign testcases[954] = 44'h92960122634;
assign testcases[955] = 44'h53881221816;
assign testcases[956] = 44'h73770131836;
assign testcases[957] = 44'h72773221837;
assign testcases[958] = 44'h74962532253;
assign testcases[959] = 44'h43891221155;
assign testcases[960] = 44'h75562411446;
assign testcases[961] = 44'h23771121254;
assign testcases[962] = 44'h33881131053;
assign testcases[963] = 44'h73561421626;
assign testcases[964] = 44'h75562411446;
assign testcases[965] = 44'h65862512625;
assign testcases[966] = 44'h92570122736;
assign testcases[967] = 44'h21596521366;
assign testcases[968] = 44'h93652612736;
assign testcases[969] = 44'h43981122153;
assign testcases[970] = 44'h65780111828;
assign testcases[971] = 44'h65780111828;
assign testcases[972] = 44'h83670122838;
assign testcases[973] = 44'h63a70121726;
assign testcases[974] = 44'h93780125726;
assign testcases[975] = 44'h22984821534;
assign testcases[976] = 44'h22984821534;
assign testcases[977] = 44'h22596732555;
assign testcases[978] = 44'h72751213533;
assign testcases[979] = 44'h5358002184b;
assign testcases[980] = 44'h54791211546;
assign testcases[981] = 44'h43681321487;
assign testcases[982] = 44'hb5854b21544;
assign testcases[983] = 44'h54791211546;
assign testcases[984] = 44'h5358002184b;
assign testcases[985] = 44'h72970111054;
assign testcases[986] = 44'h72650011627;
assign testcases[987] = 44'h22984821534;
assign testcases[988] = 44'h22571421234;
assign testcases[989] = 44'h62561321627;
assign testcases[990] = 44'h22571421234;
assign testcases[991] = 44'h21984721424;
assign testcases[992] = 44'h21862721233;
assign testcases[993] = 44'h21984721424;
assign testcases[994] = 44'h215b5422738;
assign testcases[995] = 44'h43882421154;
assign testcases[996] = 44'hb3c40021061;
assign testcases[997] = 44'hb3c40021061;
assign testcases[998] = 44'h21560111586;
assign testcases[999] = 44'hb2920111063;



winered_tnn1_tnnpar dut (.features(features),.prediction(prediction));

integer i,j;
initial begin
    features = testcases[0];
    for(i=0;i<TEST_CNT;i=i+1) begin
        features = testcases[i];
        #period
        for(j=0;j<CLASS_CNT;j=j+1) begin
            $write("%d ,",dut.scores[j]);
        end
        $display("");
    end
end

endmodule
