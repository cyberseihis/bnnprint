module tbtseqq ();

parameter N = 11;
parameter M = 40;
parameter B = 4;
parameter C = 7;
parameter Ts = 5;


parameter Wvals = 440'b00010001000000000100111010000100000100000000001110011010101111111000000011011110011000101001111010100011100000001001001001001010001000101010000001010010101000001100001001010100100000010001001010100000000110000010100011001001000001110110000101000110111100011011000110010000000101011100001001001000101001010000001111000000001000000001010000000111000000000001000001101000000000101000000000010010000110000110100001000000100010110100010100000001;
parameter Wzero = 440'b10011001110000000100111010000101000100011001101110011010111111111100011111111110011001101001111010110011101101001011101001001110011000111011011011110110101101001111101101010110110110010101001010110101001110011011110011011011100001110110110101110111111100111011101110010000001111011111011101101011111011011100011111011001101000001101010101100111000001000001000111101010100110101001010000010110000111000110100101011110101011111110110100000011;
assign data = 44'h53352264442;
parameter Wnnz = 320'h06070806070407070707040806050804090607070707080808050305010906050503060906060307;

  wire [B*N-1:0] data;
  wire [M-1:0] bitz;
  wire done;
  reg rst;
  reg clk;

  /* assign data = 16'h1234; */
  

  // Instantiate module under test
 tseqq #(
  .N(N),
  .B(B),
  .M(M),
  .Wvals(Wvals),
  .Wzero(Wzero),
  .Wnnz(Wnnz)
 ) dut (
    .data(data),
    .clk(clk),
    .rst(rst),
    .done(done),
    .out(bitz)
  );
  
  always #5 clk <= ~clk;

  integer i;
  initial begin
    /* $monitor("sums %h %0t",dut.sums,$time); */
    /* $monitor("1done %h %0t",dut.layers.layer1.done,$time); */
    runtestcase();
    $finish;
  end

  task runtestcase(); begin
    rst <= 1;
    clk <= 0;
    #10
    rst <= 0;
    #10
    #((N-1)*10)
    $display("DONE");
    $displayb(bitz);
  end
  endtask

endmodule
