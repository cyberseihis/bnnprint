












module Har_bs #(

parameter N = 12,
parameter M = 40,
parameter B = 4,
parameter C = 6,
parameter Ts = 5


  ) (
  input clk,
  input rst,
  input [N*B-1:0] data,
  output [$clog2(C)-1:0] klass
  );

  localparam Weights0 = 480'b111010100100110001110010001111111101001100000101000001000110101011100001001011000011100101111101101010010110010111000010101000001001010101010101111001000010001110000011110010011010001110100000010111011101001010000101111011111010010001111110010000001110001011011110110000000111110100000100100110101110111001001100110010010000110001101100101110000101111110000010111011111001000101010101100001000011101001100011111100011000010010100010010101011100001111100001000011010111011010111100 ;
  localparam Weights1 = 240'b001000111100001110010000101000100100111010000011111100011000110000000110111111101011001011010011101101010110011000101010010101000100001110101100011110111110011100101110010110101010010100111111011010110001010001101001111101000001101111100111 ;

  localparam SumL = $clog2(M+1);
  wire [SumL*C-1:0] sums;

  seqlego #(.N(N),.B(B),.M(M),.C(C),.Weights0(Weights0),.Weights1(Weights1)) layers (
    .clk(clk),
    .rst(rst),
    .data(data),
    .out(sums)
  );

  argmax #(.N(C),.I($clog2(C)),.K(SumL)) result (
     .inx(sums),
     .outimax(klass)
  );

endmodule
