











module cardio_tnn1_tnnseq #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnn #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(760'b1110100010000000000010000001001010000001000110000001000001000000001000010111101000000000000001010000010000010000000001100100100100010100101000000010000000000000010001111000100000100101001000000001000100000010001000000001000000100001100000001000000010001000001000011000010000100010000000101100010010010000000010000000000000000000000010010000010011000000000100000100000011001000001010000001111011101000100100001100101000011010010010000000110010110001100000010001000001000100000000001100000001000000000000010001100001100000110101111001100000010111000000000000000100000000100000000000100000001110101001010011000101000111001001100010000000000100000000000100000000011000000100000001001100110101110111010101011000100000000001011000111000000001000000000000001010111100),
  .MASK(760'b1110101110100110000010000011011110000001111110101111000001001001001000010111101101001000101001010010110000010000010101100100100111110100101000001011110011111000110001111011100010110101001010110101010100000110111010000001100000100001100110101000101010101011001000111000010010110110000010101100010010010001100011000010010000110000100011110001110011100101100100000111001111011101001110111011111111101000100100001100101010011110110011100011110011110101100011010101101111000110100010101100000101000001000111110111100101100000110111111001100011110111100000100010101100110010111110001000100000101110101101011111010111000111001011111011011011101100001010111100000010011000101100000001011111110111110111010111111110111110111111111000111001110011101000000010001011111100),
  .NONZERO_CNT(640'h0b0b090909070c0a110c09080a0906090804090b0d08080a0b040d08080b0a070b090c0c0a0a0807),
  .SPARSE_VALS2(39'b101110010111100011111111011101111110001),  // Bits of not-zeroes
  .COL_INDICES(312'h26211f1b130f0d0b080705040225211e1c1b0f0c090706050201252421201c1b1a18110c0a0301), // Column of non-zeros
  .ROW_PTRS(32'h271a0d00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
