












module pendigits_bnn1_bnnshift #(

parameter FEAT_CNT = 16,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 10,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 640'b0111100101011001111011000111010001000000100011110110010000110111100011000011011001110011010010011110010001111000010000011110110000011010110111100101000000001100100010100110110100110101000111000011001101010000000111110111000000100010110010101100101010100111101111011001111000111001001101101111100101110100100000101101011101011111001000111011010010010000000111001101111111010000100101101001100000111101100011100010101110001000111100011011110001001111110101111000111100101100110101100101001101010110010010111100011111011010001010000010001010101000101101010100100010100001110011000000000101101011011000111110100000001111111110110111111100001000 ;
  localparam Weights1 = 400'b0000100000101111101101100001011000110000011110110111101011101100111100000000000001011101010001011000011110000100011101100111000000001111010000000110111100001000010010110010110110100000011111111101000010001000011011000111010110000010000010110101011011010111100111100010101011111110110001011100011000001010100011000011111010001111111000101011111010000101001111000111000011011001011111000001101001000001 ;

  seq_bnn #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
