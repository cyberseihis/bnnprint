












module cardio_bnn1_bnnseq #(

parameter FEAT_CNT = 19,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 3,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 760'b0011100010010101010110101000111001101000011010010101000110110011100000010001101101001011111100011010011110011001101101010100110000010010011101010100000110000011000001011110100001000100010000100101111111001010001010010100110111001001001100101001100110001010001011000100101111001101011001110000010100001110000010000101100010101001100111011010001101001101000110101011000000000111110000000010101001001100110000011011110000100010011111111111000110100101110110110011101011011001100100111010110011101110001000000010001010000100101110010010110110000111001001011101101100010011000101101000010010111010011111000110100110111000001001110101000110110011101001101001010001001001101100101010000001000001101110010010011101010001000100110000110100101010100110001100111101101101 ;
  localparam Weights1 = 120'b101010000001111100000011001000100011100111001011000110110011011101101001101001110100101100111001001101110110000110110011 ;

  seq_bnn #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
