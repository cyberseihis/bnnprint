











module Har_ts #(

parameter FEAT_CNT = 12,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnn #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(480'b000001000100011011010000000001110000000111000001010001010000000001010001111110000001011100010010000000010010000010000000010110100011000110100000110101110000100100000000000010000000100001000100011100100100010011001000001100100000100000000000100011010000101000010100111001000100010000001100000111100000010110001000011001011100110100100000110110000000001100000010010001100110100000101000110100000001000010000000000001100001001100100000001100011000001101001000001110011000000000100000),
  .MASK(480'b100101010100111111110001010011110111111111000011111001010101100011110111111110000101011111110010000100010110011011000100110110111111011110110100111101111110100110110001001010000000101101110101111110110101010111101101001100100000100111001100100011010100101001010100111101010111010011001101010111100001011111101101011001011100111100100000111110101000101100010011110111110110110011101111110110101001010110001000110101111001101100100000101110011011101101011101111110011100110011110011),
  .NONZERO_CNT(640'h0a0702070707060b050a0705070806060606060a0604060707090705060806080809080806060408),
  .SPARSE_VALS2(89'b10010110011111001000011111001110110110101011011001101110001000101101101100100001101100111),  // Bits of not-zeroes
  .COL_INDICES(712'h272623201d1b1a1712110d0b03002623201f1d19120e0c0b0805042622201f1d18151211100b04010021201b1a1918161512110d0a060100242322211f1d18161412100e0c0b0a06052422201e1c1a1918161411100e0d0a06), // Column of non-zeros
  .ROW_PTRS(56'h594b3e30211000) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
