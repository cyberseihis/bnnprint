
















module winewhite_bnn1_bnnpaarter #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1000


)(
    input [FEAT_CNT*FEAT_BITS-1:0] features,
    output [$clog2(CLASS_CNT)-1:0] prediction
);

localparam PAAR0 = 4752'h001600530001001b005200010007005000010010004e0001001500470001001800450001001f00430001001500420001001600390001002000380001001c00320001002a00310001001f002e00010026002a0001001d00290001002100250001001600220001001600210001003400480000003500460000002d00440000001b003c00000028003b00000027003a0000001d00370000002300360000002000330000001300310000001a002e00000026002d00000019002c00000011002c0000001c002b00000016002b0000001d002a0000001a00290000001600290000001f00280000001a00280000001700260000001100250000000700250000001e00240000001d00240000001f00220000001c00220000001a00220000001c00210000001a002100000013001d00000015001c00000013001c0000000d001b00000010001a0000000f001800000016001700000011001500000007001300000007000b00000015002400000012001400010016002f0000000d00270000000b00230000001700200000001300160000001100180000000d001b0001000d00190001000f00170001000f00100001001200140000000e001400000011001700010011001e0000001300190001000f00180001000f00130000000c001200000007000d0000000e00140001000c000e0001001000110000000c00120001000f00100000000b00150001000100030000000c000e00000007000d00010005000600000000000400010002000900010008000a00000007000b00010008000a0001000200090000000000040000000500060001000100030001 ;
localparam YMAP = 1280'h0000004c0000006800010067000000620001004f0000005d0000003d000000600000006b0001005100010061000100410000004b000000490000004d0000005a00010056000000690001003f000000300001005f0001005400010055000100590001005c000100580000006d0000006400000040000100630000003e000100660000004a0000005e00000030000100650000005b0001006c000100570001006a;
localparam ADDCNT = $bits(PAAR0) / 48;
localparam FULLCNT = ADDCNT + FEAT_CNT;
localparam Weights1 = 280'b1100111000000011001100101100101011000111100011011110001100111111010011101101011100011011111010110001111101001110110101110000110111101010000011000100001011010011000011011110101100001111010011101101011100001101100010110001111111101110111001110000000011001010100110110101111011010110 ;
localparam WIDTH = 320'h07070606060706070707070606060707060606060708060706060606060706070706060607060707;
localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
localparam INDEX_BITS = $clog2(FEAT_CNT+1)+FEAT_BITS;
wire signed [FEAT_BITS:0] feature_array [FEAT_CNT-1:0];
wire [HIDDEN_CNT-1:0] hidden;
wire [HIDDEN_CNT-1:0] hidden_n;
wire [CLASS_CNT*SUM_BITS-1:0] scores; 
assign hidden_n = ~hidden;

wire signed [INDEX_BITS:0] node [FULLCNT-1:0];

genvar i;
generate
    for(i=0;i<FEAT_CNT;i=i+1)
        assign feature_array[i] = {1'b0,features[i*FEAT_BITS+:FEAT_BITS]};
    for(i=0;i<FEAT_CNT;i=i+1)
        assign node[i] = feature_array[i];
endgenerate

integer j;
generate
for(i=0;i<ADDCNT;i=i+1) begin
    localparam adsub = PAAR0[i*48];
    localparam op1 = PAAR0[i*48+16+:16];
    localparam op2 = PAAR0[i*48+32+:16];
    localparam nodeloc = FEAT_CNT + i;
    if(adsub)
        assign node[nodeloc] = node[op1] + node[op2];
    else
        assign node[nodeloc] = node[op1] - node[op2];
end
for(i=0;i<HIDDEN_CNT;i=i+1) begin
    localparam ymap = YMAP[i*32+:16];
    localparam signy = YMAP[i*32+16];
    if(signy)
        assign hidden[i] = node[ymap] >= 0;
    else
        assign hidden[i] = node[ymap] < 0;
end
endgenerate

initial begin
    #10
    for(j=0;j<FULLCNT;j=j+1) begin
        $display("%d | %d | %b, %d, %d", j, node[j], PAAR0[(j- FEAT_CNT )*48],  PAAR0[(j-FEAT_CNT)*48+16+:16], PAAR0[(j-FEAT_CNT)*48+32+:16]);
    end
end

generate
for(i=0;i<CLASS_CNT;i=i+1) begin
    localparam Wneur = Weights1[i*HIDDEN_CNT+:HIDDEN_CNT];
    reg unsigned [SUM_BITS-1:0] tmpscore;
    always @ (*) begin
        tmpscore = 0;
        for(j=0;j<HIDDEN_CNT;j=j+1) begin
        if(Wneur[j])
            tmpscore = tmpscore + hidden[j];
        else 
            tmpscore = tmpscore + hidden_n[j];
        end
    end
    assign scores[i*SUM_BITS+:SUM_BITS] = tmpscore;
end
endgenerate

argmax #(.SIZE(CLASS_CNT),.INDEX_BITS($clog2(CLASS_CNT)),.BITS(SUM_BITS)) result (
    .inx(scores),
    .outimax(prediction)
);
endmodule
