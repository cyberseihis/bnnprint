`timescale 1us/1ns





module tbpendigits_ts #(

parameter FEAT_CNT = 16,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 10,
parameter TEST_CNT = 1000




)();
  reg [FEAT_BITS*FEAT_CNT-1:0] data;
  wire [FEAT_BITS*FEAT_CNT-1:0] testcases [TEST_CNT-1:0];
  reg rst;
  reg clk;
  parameter Nsperiod=50000;
  localparam period=Nsperiod/500;
  localparam halfT=period/2;


assign testcases[0] = 64'h8f4d96400498fe6f;
assign testcases[1] = 64'h0e4f7c572260b0f1;
assign testcases[2] = 64'h095bceffcc884430;
assign testcases[3] = 64'h0f1f1b37e5f7c4b0;
assign testcases[4] = 64'h0b8dffddaa665380;
assign testcases[5] = 64'hffef8c380360c333;
assign testcases[6] = 64'h0f0c46e6fbcfa8b0;
assign testcases[7] = 64'h060a21a0f7ef6f09;
assign testcases[8] = 64'h2e28c690130a5fff;
assign testcases[9] = 64'h9f4c0540c2f8ce4e;
assign testcases[10] = 64'hce5f0baafdf6d030;
assign testcases[11] = 64'h8faae43035dbff0e;
assign testcases[12] = 64'hffcf6c59d8a23000;
assign testcases[13] = 64'hfc9f0e49dbf6d130;
assign testcases[14] = 64'h0e6fdee8d29084f4;
assign testcases[15] = 64'h6c9fffbbd6d15003;
assign testcases[16] = 64'h8dbfcc88f7f28001;
assign testcases[17] = 64'hfdaf4cdbfaf49003;
assign testcases[18] = 64'h4b7f9a54003290f0;
assign testcases[19] = 64'h0c3fcfbc581370f0;
assign testcases[20] = 64'h2c3ac680030a4fff;
assign testcases[21] = 64'h078acefffce8c4e0;
assign testcases[22] = 64'h2e5bb550140b5fff;
assign testcases[23] = 64'hca8f0cd6f02289ef;
assign testcases[24] = 64'h9f5c1702b0f47763;
assign testcases[25] = 64'h2f0b27e8facbb5b0;
assign testcases[26] = 64'h6f1d0640c1f7de6f;
assign testcases[27] = 64'h7f2d5afcbd894400;
assign testcases[28] = 64'ha99f0d77d01157fb;
assign testcases[29] = 64'hfd5f0e1b28260300;
assign testcases[30] = 64'h598fffd780f3990a;
assign testcases[31] = 64'h6f8bd460041c7fff;
assign testcases[32] = 64'h0f6fdeb7904486f5;
assign testcases[33] = 64'h4c0730b0f6fd7f0c;
assign testcases[34] = 64'h0052a5e8fddf9dda;
assign testcases[35] = 64'h5ebfcc88c6f39001;
assign testcases[36] = 64'h5f29b650030c6fff;
assign testcases[37] = 64'hcf6f0915d5fac780;
assign testcases[38] = 64'haf0bfbef2bfbf640;
assign testcases[39] = 64'h1f8fed98350180f0;
assign testcases[40] = 64'h0faffcb7816026e6;
assign testcases[41] = 64'h5e39b780032a7fff;
assign testcases[42] = 64'haf3c0620b0f59622;
assign testcases[43] = 64'h0d5fefabc7f28020;
assign testcases[44] = 64'h1e7feffdc9a56200;
assign testcases[45] = 64'hffbf4b0540f1c619;
assign testcases[46] = 64'h8ecfecb8f4d16002;
assign testcases[47] = 64'h5c7fcca7420181f0;
assign testcases[48] = 64'h0e099560241b4fff;
assign testcases[49] = 64'haf6cbafcdc985400;
assign testcases[50] = 64'h2f9fdd89e6f29000;
assign testcases[51] = 64'h8cbfffdd9a562300;
assign testcases[52] = 64'h9f3c0460e4fb9f3c;
assign testcases[53] = 64'h0c8efffdca866330;
assign testcases[54] = 64'h3f0c16c6facfb8c0;
assign testcases[55] = 64'h7f3c8650050e8fff;
assign testcases[56] = 64'h3daffdb9d8e37002;
assign testcases[57] = 64'h2c6fcc87220381f0;
assign testcases[58] = 64'h3c0c2490f4fb8f1d;
assign testcases[59] = 64'hff7e190480f48612;
assign testcases[60] = 64'h9aff0f68f30016fb;
assign testcases[61] = 64'h5defff6e79f59000;
assign testcases[62] = 64'h2a0370f4fabf2f08;
assign testcases[63] = 64'h0d8fcd6887f4a000;
assign testcases[64] = 64'h0fafffaa65201587;
assign testcases[65] = 64'hfdbf4c76800166f9;
assign testcases[66] = 64'h6fdfff8e59c67000;
assign testcases[67] = 64'hff9d593470d38706;
assign testcases[68] = 64'hfd6f2a95b00378fd;
assign testcases[69] = 64'h0dc9f24047fcdf0d;
assign testcases[70] = 64'hdf6f9dadd8f28001;
assign testcases[71] = 64'h6c0720a1f7fe8f1b;
assign testcases[72] = 64'h5f3c0675f5f7c7b0;
assign testcases[73] = 64'h0c5cbdfffdd9b490;
assign testcases[74] = 64'hebff4e28daf8a300;
assign testcases[75] = 64'h0f7fbb86503467f7;
assign testcases[76] = 64'h6f1a0370d3facf5f;
assign testcases[77] = 64'hcf6e090380f39521;
assign testcases[78] = 64'h4dbffe99e7f28000;
assign testcases[79] = 64'h1c8fffbbf7f27002;
assign testcases[80] = 64'h5c9f98520052a0f0;
assign testcases[81] = 64'h7f3e0a47b7f8c490;
assign testcases[82] = 64'h7bcfcd96700281f2;
assign testcases[83] = 64'h5f2c080360f1a330;
assign testcases[84] = 64'h3e1a8640160d8fff;
assign testcases[85] = 64'h3e09e9e320172dff;
assign testcases[86] = 64'h0f9ffeb8a3c0f576;
assign testcases[87] = 64'h8f0b0380f5fd7f1a;
assign testcases[88] = 64'h681b0370e4fbaf3d;
assign testcases[89] = 64'hff8f3ccefeb96400;
assign testcases[90] = 64'h3e096400053b7fff;
assign testcases[91] = 64'h6f4d080380f3b719;
assign testcases[92] = 64'h4f0b0585f6dac5b0;
assign testcases[93] = 64'h0f8fdbd4c0f58707;
assign testcases[94] = 64'h0a6dafcecad7d3f0;
assign testcases[95] = 64'h3d072090e5fbcf5f;
assign testcases[96] = 64'h0a6ddfffdba79490;
assign testcases[97] = 64'h6c38fbbf0ca9f8f0;
assign testcases[98] = 64'hffac480410a0c443;
assign testcases[99] = 64'h593ecffa840060f0;
assign testcases[100] = 64'h2f1842c0f6ed7f0d;
assign testcases[101] = 64'h3eafbc78f8f38000;
assign testcases[102] = 64'h1f0b34a0f3fa9f1c;
assign testcases[103] = 64'h7da8e22005c9ff3f;
assign testcases[104] = 64'h1a2280f2facf4f0a;
assign testcases[105] = 64'h6feffd99b5f29000;
assign testcases[106] = 64'h492a0370e4fbbf5b;
assign testcases[107] = 64'h4f0921a0f6ff8f38;
assign testcases[108] = 64'h7f2b8630160d7fff;
assign testcases[109] = 64'h0e6f3b17e8f9d4e0;
assign testcases[110] = 64'hcf6f0902b1f75710;
assign testcases[111] = 64'h2c0550d0f6ec7f3b;
assign testcases[112] = 64'hef5d190480f3b806;
assign testcases[113] = 64'h0e4bc57055dbff1e;
assign testcases[114] = 64'h8fcbff7efce8b100;
assign testcases[115] = 64'h7f1d0785f7e87530;
assign testcases[116] = 64'h1f098660121a7fff;
assign testcases[117] = 64'hfcff8c380260c454;
assign testcases[118] = 64'h7bbfda84100081f1;
assign testcases[119] = 64'h6f89cf4fdbf48004;
assign testcases[120] = 64'hfe6da6d00188df0c;
assign testcases[121] = 64'h7f0acbe530274fff;
assign testcases[122] = 64'h7f2b1390f5fd6f0a;
assign testcases[123] = 64'h2b2570e3f9de5f0c;
assign testcases[124] = 64'h8d190380f4fbaf1e;
assign testcases[125] = 64'h3f0c1975f6f8f4e0;
assign testcases[126] = 64'h4f0f8fffbd794450;
assign testcases[127] = 64'h8fcfeb97f7e27002;
assign testcases[128] = 64'hff8f8cfffeb96400;
assign testcases[129] = 64'h5c9fbb76220181f0;
assign testcases[130] = 64'h2f1a7660240c8fff;
assign testcases[131] = 64'h8e58fabf9bfab000;
assign testcases[132] = 64'hbf4d0720a0f5fb9e;
assign testcases[133] = 64'hffaf5c2711707405;
assign testcases[134] = 64'hfb9f2c0480f3fb7d;
assign testcases[135] = 64'hdf9f3c0732f0f414;
assign testcases[136] = 64'hff8d492460f1a504;
assign testcases[137] = 64'h07599cefffdba680;
assign testcases[138] = 64'hbf5e0976f8fbb560;
assign testcases[139] = 64'hce5a0081f9dfdc64;
assign testcases[140] = 64'h4d0650d1f9bf4f18;
assign testcases[141] = 64'hef8d280470f3c616;
assign testcases[142] = 64'h6dafcc770301a0f0;
assign testcases[143] = 64'hfebf3dbefbb76300;
assign testcases[144] = 64'h5f3a8470250b4fff;
assign testcases[145] = 64'h0c7fffccf6f07004;
assign testcases[146] = 64'h0759adfffed9a470;
assign testcases[147] = 64'h3f1c0876f8f8e4c0;
assign testcases[148] = 64'h0b3f4b250051b2f2;
assign testcases[149] = 64'h8f6d380383f5f6f0;
assign testcases[150] = 64'h56aafdffcc884400;
assign testcases[151] = 64'h0a7cdfffecc8b4d0;
assign testcases[152] = 64'h088dfff9d23031f1;
assign testcases[153] = 64'haf4d0812a0f49807;
assign testcases[154] = 64'hed2dffffab571400;
assign testcases[155] = 64'h2d8bff4f0bdcc680;
assign testcases[156] = 64'h0d89f580448acf1f;
assign testcases[157] = 64'hcf6d2a0664e5f4d0;
assign testcases[158] = 64'h0fbfec96501557f7;
assign testcases[159] = 64'h6dbffe9ae6f18000;
assign testcases[160] = 64'h0fcffdfaf8d5a240;
assign testcases[161] = 64'h09ccff3f1bdb7630;
assign testcases[162] = 64'h0e5fcca680f1b507;
assign testcases[163] = 64'h2f0c48f9fcfbf5f0;
assign testcases[164] = 64'h3c6fefbaf7f28002;
assign testcases[165] = 64'h8f2d0640b0f5ec7f;
assign testcases[166] = 64'h4ffffca8633005c6;
assign testcases[167] = 64'h7effff8e1a888300;
assign testcases[168] = 64'h9f0e97b01198ff1f;
assign testcases[169] = 64'h7deffdc9e6f28002;
assign testcases[170] = 64'hdf7f2a0380f55621;
assign testcases[171] = 64'h4c38a330040a7eff;
assign testcases[172] = 64'h6acedf9a650051f0;
assign testcases[173] = 64'h2f098860021b7fff;
assign testcases[174] = 64'h0a7cffffbc884410;
assign testcases[175] = 64'h0b8eafacb9d6f2f0;
assign testcases[176] = 64'h0b3dafefece8f4f0;
assign testcases[177] = 64'hef7dcceffbf69100;
assign testcases[178] = 64'h5f3d0844d5fad5b0;
assign testcases[179] = 64'h4f29c89010096fff;
assign testcases[180] = 64'h0c3f9fffedb98580;
assign testcases[181] = 64'h0f7fedf6e0f4f888;
assign testcases[182] = 64'h3fefebb5800447f7;
assign testcases[183] = 64'h5f1a0450c3f8de6f;
assign testcases[184] = 64'h3c9ffffce8c47100;
assign testcases[185] = 64'hff8c380440f1f544;
assign testcases[186] = 64'hdc3b2fbffcc76300;
assign testcases[187] = 64'hff9d490400909303;
assign testcases[188] = 64'h3e6cff0facf8b440;
assign testcases[189] = 64'h390550c2f9ef6f1b;
assign testcases[190] = 64'hde7f0c9bffeac5c0;
assign testcases[191] = 64'h0f7f9a73401695f5;
assign testcases[192] = 64'h0badeffefbf7d4b0;
assign testcases[193] = 64'h5f1b0450b2f7fdaf;
assign testcases[194] = 64'hffbf7d89f8d37000;
assign testcases[195] = 64'h8f3b0530b1f5fc8e;
assign testcases[196] = 64'hffaf4e6ac9c47000;
assign testcases[197] = 64'h589bffedc8b300f1;
assign testcases[198] = 64'hee6f3cdcfcf5a001;
assign testcases[199] = 64'hbf6d0a16b6f8c490;
assign testcases[200] = 64'h8f4c09cbfdbe7730;
assign testcases[201] = 64'h4f0c69f9df9a7550;
assign testcases[202] = 64'h0d689210071c8fff;
assign testcases[203] = 64'h8ffffcc8740170f0;
assign testcases[204] = 64'hffbf6b2702608404;
assign testcases[205] = 64'h9f0e78f3a0a6ed4f;
assign testcases[206] = 64'h0a4e9fcc875290f1;
assign testcases[207] = 64'h0c5dbfffdcb89390;
assign testcases[208] = 64'h084aadfffde9c4a0;
assign testcases[209] = 64'h6eefec88f7f38000;
assign testcases[210] = 64'hceabf480259bbf0d;
assign testcases[211] = 64'hbf5c69eafda95400;
assign testcases[212] = 64'h0e9ffdc7803255f6;
assign testcases[213] = 64'hfffecb9997541200;
assign testcases[214] = 64'h8f6aa430160f8fff;
assign testcases[215] = 64'h0f7fffddaa776350;
assign testcases[216] = 64'h2c5ab550150b6fff;
assign testcases[217] = 64'hdf3f48700499ff4f;
assign testcases[218] = 64'h6d3a6320053c8fff;
assign testcases[219] = 64'h8f5c0837b6f9e5e0;
assign testcases[220] = 64'hcf6f391380f46500;
assign testcases[221] = 64'h0e8feeca762270f0;
assign testcases[222] = 64'h7ddffec9f6f28000;
assign testcases[223] = 64'hdfac480472f5f4f0;
assign testcases[224] = 64'h8f0e19fafbedb6e0;
assign testcases[225] = 64'hfbcf3ca6b00258fd;
assign testcases[226] = 64'hffbe592480f3b708;
assign testcases[227] = 64'h5a8f99630043a0f1;
assign testcases[228] = 64'h6f2c7740011a6fff;
assign testcases[229] = 64'h4f489430052e8fff;
assign testcases[230] = 64'hff8d381370f29504;
assign testcases[231] = 64'h0f6fab94703697f7;
assign testcases[232] = 64'h0d4f8c75500585f6;
assign testcases[233] = 64'h085baeffdca88450;
assign testcases[234] = 64'h0f8fffca957035b6;
assign testcases[235] = 64'h296a9f9a93f28100;
assign testcases[236] = 64'h7fdfdccaf6c26001;
assign testcases[237] = 64'h0b6ba560157afe9f;
assign testcases[238] = 64'hfc5a0e8ffdf8a430;
assign testcases[239] = 64'h5c0710a0f5fc8f0d;
assign testcases[240] = 64'h8ddffc98f8e27003;
assign testcases[241] = 64'h5f190360c3f9ff8f;
assign testcases[242] = 64'h0f7fcc96604487f6;
assign testcases[243] = 64'hfcff4d67b10075fa;
assign testcases[244] = 64'h1a4f9c74011483f0;
assign testcases[245] = 64'hafdbff6fbaf7a100;
assign testcases[246] = 64'hcf8e0720e5fdc821;
assign testcases[247] = 64'h0062b5fafeaf7cc8;
assign testcases[248] = 64'h89fcaf0d2aeaf5e0;
assign testcases[249] = 64'h070a8dfffcc87450;
assign testcases[250] = 64'hcf7b0747f7eaa590;
assign testcases[251] = 64'hffbf5a0450d39808;
assign testcases[252] = 64'h0d6fdd7897f4a001;
assign testcases[253] = 64'h0c4fbfda944090f0;
assign testcases[254] = 64'hffbc692520807303;
assign testcases[255] = 64'h4f0c1390f6de5f37;
assign testcases[256] = 64'hff2ec9df6a066067;
assign testcases[257] = 64'hbf3c0550d5fc9f2c;
assign testcases[258] = 64'hef0f59f45016db8f;
assign testcases[259] = 64'hcd5c0d9ffec86400;
assign testcases[260] = 64'h5dbfdc88f8f27002;
assign testcases[261] = 64'h0bc7f13066fcef1d;
assign testcases[262] = 64'hffaf6c3823406406;
assign testcases[263] = 64'hef9c7691f0f57604;
assign testcases[264] = 64'h4c9ffdb8540081f3;
assign testcases[265] = 64'h5e181190f5fb9f0f;
assign testcases[266] = 64'ha7fcbf1e09c9f5f0;
assign testcases[267] = 64'h0e7fefffdcb894a0;
assign testcases[268] = 64'h6c1a0280f5fd8f3a;
assign testcases[269] = 64'h9d4ae44046fccf0c;
assign testcases[270] = 64'hce0f3ad5b0145aff;
assign testcases[271] = 64'h0f1d0925a4f7f4e0;
assign testcases[272] = 64'hbf7b260485f7f6e0;
assign testcases[273] = 64'haf4f0923a0f38410;
assign testcases[274] = 64'hff8f3b0540d1d554;
assign testcases[275] = 64'h2f1f0b1796f8d4b0;
assign testcases[276] = 64'h2f0840c0f7de5f0a;
assign testcases[277] = 64'h49acffcb97620040;
assign testcases[278] = 64'h7d8fdfb8730081f0;
assign testcases[279] = 64'h0d5fcdd7c16073f3;
assign testcases[280] = 64'h5d4feffbd7f37004;
assign testcases[281] = 64'h7f0b04b4f8cfd8e0;
assign testcases[282] = 64'hffbfaeeec8b36002;
assign testcases[283] = 64'hffad694470d27403;
assign testcases[284] = 64'hff9f4d3888b46001;
assign testcases[285] = 64'h6b5fae78031390f3;
assign testcases[286] = 64'hff9c480430d1b514;
assign testcases[287] = 64'h0f8ffdd7b17005d6;
assign testcases[288] = 64'hffae592530f1b402;
assign testcases[289] = 64'hff6f2d46c8f39001;
assign testcases[290] = 64'h4c8fffdba8d38001;
assign testcases[291] = 64'h4b7fcd88230080f1;
assign testcases[292] = 64'hffaf3c27b8e37001;
assign testcases[293] = 64'hff9e3b0631b0b548;
assign testcases[294] = 64'hcf5c0898fcc98460;
assign testcases[295] = 64'h6dcffcb8f7f38000;
assign testcases[296] = 64'h78affeb750c39a0c;
assign testcases[297] = 64'h0d5fbea75343a2f0;
assign testcases[298] = 64'h5e49c68002297fff;
assign testcases[299] = 64'h2d8fffdbc8e37002;
assign testcases[300] = 64'h9effff8e4aa58000;
assign testcases[301] = 64'h0f7fffda853035c6;
assign testcases[302] = 64'h8f3d0936a6f7d4a0;
assign testcases[303] = 64'h2c7ffeb9c8f28003;
assign testcases[304] = 64'hff9f4d6bc9c47000;
assign testcases[305] = 64'h0559acffece8d4d0;
assign testcases[306] = 64'h0c4fcffde99561d0;
assign testcases[307] = 64'hffbf5e4999a46000;
assign testcases[308] = 64'hfa8f0d87e17097fd;
assign testcases[309] = 64'h15aadf1f69f49004;
assign testcases[310] = 64'h7f5c0707a6f9f6e0;
assign testcases[311] = 64'h0c6ffcb670f1664c;
assign testcases[312] = 64'h7fffcf6ba8f38002;
assign testcases[313] = 64'hfc7a0c6fced9c4e0;
assign testcases[314] = 64'h5cbffeaaf7d27001;
assign testcases[315] = 64'h2e0750d1faaf4c53;
assign testcases[316] = 64'h0e5fcfba672381f0;
assign testcases[317] = 64'h0d6fcba5501477f7;
assign testcases[318] = 64'h3d299f4e666001f1;
assign testcases[319] = 64'h0a7f8f8a841021f0;
assign testcases[320] = 64'h6a0b8dffdcb88380;
assign testcases[321] = 64'h2f4f0a06b6f9d5b0;
assign testcases[322] = 64'h0e7fcda6806287f7;
assign testcases[323] = 64'h0e7feffad5a04395;
assign testcases[324] = 64'h9c4bb56085fbbf0e;
assign testcases[325] = 64'h086ccfffcc886440;
assign testcases[326] = 64'h7f3f7b9febf49000;
assign testcases[327] = 64'h4f0921a0f5fd7f0c;
assign testcases[328] = 64'hffbf4b0620c0c528;
assign testcases[329] = 64'h6c9f3a0470f47641;
assign testcases[330] = 64'h4bfe5be55005accf;
assign testcases[331] = 64'h6f9f88430353b1f0;
assign testcases[332] = 64'h1e8fdc98e7f49000;
assign testcases[333] = 64'hff1f7ae5900268fc;
assign testcases[334] = 64'h0e4fae7a1743a2f0;
assign testcases[335] = 64'h7f1bcca400183fff;
assign testcases[336] = 64'h4daffc8896f39001;
assign testcases[337] = 64'hff7f1a0470f47530;
assign testcases[338] = 64'h0d6fdeaaf7f29021;
assign testcases[339] = 64'h0c4fafaa651180f0;
assign testcases[340] = 64'h0f6f9ca8744190f0;
assign testcases[341] = 64'hff9c482450e1a403;
assign testcases[342] = 64'h1d3f4b250050b1f1;
assign testcases[343] = 64'h8e3a0430b1f6fbaf;
assign testcases[344] = 64'hed8f3aa4b00076fb;
assign testcases[345] = 64'h6f8bcf4efdf59005;
assign testcases[346] = 64'h0fafbb85502256f7;
assign testcases[347] = 64'h0b29b68022395fff;
assign testcases[348] = 64'hcf8a0697f9eca680;
assign testcases[349] = 64'h6dafed8af8f49100;
assign testcases[350] = 64'h0c7effddb99692a0;
assign testcases[351] = 64'h7a0c8fffdcc8c4f0;
assign testcases[352] = 64'hffcd793450c18404;
assign testcases[353] = 64'hff9f5aecfef8a200;
assign testcases[354] = 64'h091280e4fbcf5d17;
assign testcases[355] = 64'h3eaffdd8840130c0;
assign testcases[356] = 64'h280360d1f7cd6f0d;
assign testcases[357] = 64'h5cbffcb6130593f0;
assign testcases[358] = 64'hec8f2c36000589fe;
assign testcases[359] = 64'h4e0a10a0f7df5f16;
assign testcases[360] = 64'h2b6fab75020181f0;
assign testcases[361] = 64'hff8e390430c0b312;
assign testcases[362] = 64'hdf5d180360f1e544;
assign testcases[363] = 64'h091b7ddfffdba5b0;
assign testcases[364] = 64'h0d8fcc86403478f8;
assign testcases[365] = 64'hfbcf1f0bbcfcf6e0;
assign testcases[366] = 64'h6cafab56032292f0;
assign testcases[367] = 64'h4c7fcb94100181f0;
assign testcases[368] = 64'h2f1b0633c3f7c5c0;
assign testcases[369] = 64'h3f2ba880230c7fff;
assign testcases[370] = 64'h3d9ffeabe6f28000;
assign testcases[371] = 64'h6f0d49faafad96a0;
assign testcases[372] = 64'h0d4f8d78442090f0;
assign testcases[373] = 64'h5dbfba65011380f1;
assign testcases[374] = 64'hff4f0b7550046aef;
assign testcases[375] = 64'h3e17a860022b6fff;
assign testcases[376] = 64'h3f0740c0f8ef7f48;
assign testcases[377] = 64'hcf0f3ad5b076fbef;
assign testcases[378] = 64'h3c8fed79e9f48003;
assign testcases[379] = 64'h1e0842c0f6dd6f0b;
assign testcases[380] = 64'h0fbfda95700355f5;
assign testcases[381] = 64'h6fcfdcb9f5c16001;
assign testcases[382] = 64'h5f2c081370f2d534;
assign testcases[383] = 64'h2c6fffb8520017b9;
assign testcases[384] = 64'h9ccfaa64002190f0;
assign testcases[385] = 64'h0669bcfffcd8b4b0;
assign testcases[386] = 64'hef9e0a78f9dc8630;
assign testcases[387] = 64'h1e0a23a0f5fc8f1c;
assign testcases[388] = 64'h0f1f9ffefac78460;
assign testcases[389] = 64'h0f8fff9950b2b454;
assign testcases[390] = 64'h8f3c080370f38411;
assign testcases[391] = 64'hac5f0922b0f6ed5e;
assign testcases[392] = 64'h0d2f9f8bb7f3c030;
assign testcases[393] = 64'hfb9f4cc5a00499cc;
assign testcases[394] = 64'hff9e390440c19504;
assign testcases[395] = 64'hffae5b1702609334;
assign testcases[396] = 64'h4d082180f4facf5f;
assign testcases[397] = 64'h6cc6d02086fbcf0d;
assign testcases[398] = 64'h6dcffba6230594f0;
assign testcases[399] = 64'h4c8fcd88d7f39001;
assign testcases[400] = 64'h2eaffe9ad7f4a001;
assign testcases[401] = 64'hdf0f1ceeffdaa590;
assign testcases[402] = 64'h0e298580343b8fff;
assign testcases[403] = 64'h0b6dcfffcc884420;
assign testcases[404] = 64'hef6d0700a0f6fe7f;
assign testcases[405] = 64'haacf2f6cfef7a100;
assign testcases[406] = 64'hcf5c180380f2c635;
assign testcases[407] = 64'h6a9f9c95c0f16101;
assign testcases[408] = 64'hdf6d190460f1e543;
assign testcases[409] = 64'h7dbffc98f7f38000;
assign testcases[410] = 64'h0f8fffe9925066f6;
assign testcases[411] = 64'hcd8fa9d30045facf;
assign testcases[412] = 64'h0cafcfbcc8d480f0;
assign testcases[413] = 64'h4a5fad97420180f0;
assign testcases[414] = 64'hfddf4f0e39b6e150;
assign testcases[415] = 64'h4ceaff5ebaf9d200;
assign testcases[416] = 64'h5c8fa963003392f0;
assign testcases[417] = 64'h2c8ffffc89c58100;
assign testcases[418] = 64'h1f0c17a4f7e9b490;
assign testcases[419] = 64'h0f7ffffdcaa68390;
assign testcases[420] = 64'h0f6fbd86403487f7;
assign testcases[421] = 64'h5f2cb65035fabf0c;
assign testcases[422] = 64'h9f4c1804b4f8d4b0;
assign testcases[423] = 64'h2d7fdd98e7f28001;
assign testcases[424] = 64'h5cfcff0d09fb7610;
assign testcases[425] = 64'h0f6fce97504287f7;
assign testcases[426] = 64'haf5cf6f00066eccf;
assign testcases[427] = 64'hff8f2e1868c48000;
assign testcases[428] = 64'h1e073180d3fadf8f;
assign testcases[429] = 64'h8e8fffdbd6e16004;
assign testcases[430] = 64'h1c0560e2fabf3c35;
assign testcases[431] = 64'hcacf2e28610055f9;
assign testcases[432] = 64'h6f3d0866f7fad5e0;
assign testcases[433] = 64'h0f8fffc9937046d8;
assign testcases[434] = 64'hffac6670f0f58804;
assign testcases[435] = 64'h5f0b469200277dff;
assign testcases[436] = 64'h1d0f6d58141180f0;
assign testcases[437] = 64'h0d5fbffefac683a0;
assign testcases[438] = 64'h8f6a05e5f9ceb7a0;
assign testcases[439] = 64'hdd6f0b13a0f5ed6f;
assign testcases[440] = 64'h4eafddcaf6d27001;
assign testcases[441] = 64'h5e1922a0f5fc8f0d;
assign testcases[442] = 64'h0d4f9c86602375f5;
assign testcases[443] = 64'h7dbfcdbaf6e27002;
assign testcases[444] = 64'h2e9fdeaaf8e47100;
assign testcases[445] = 64'h2f0c57f9ffdde7f0;
assign testcases[446] = 64'h9effef8c97e48000;
assign testcases[447] = 64'h5fff9f0b17c5c120;
assign testcases[448] = 64'h0f7fddf8f2e0e474;
assign testcases[449] = 64'h0f8ffee8b28045c7;
assign testcases[450] = 64'h0f3f1a46b7f9e4f0;
assign testcases[451] = 64'hbfffdf8d88934002;
assign testcases[452] = 64'h7f1a0270d4fcaf3f;
assign testcases[453] = 64'hcf6f6ddffdb86300;
assign testcases[454] = 64'h0a6ddffeeab69280;
assign testcases[455] = 64'h6fff7f0c4ae7c330;
assign testcases[456] = 64'h5c9fcb96310180f1;
assign testcases[457] = 64'hffdd690410c1b524;
assign testcases[458] = 64'h2c8fee8ac6f18002;
assign testcases[459] = 64'h0a8dfffdaa8673a0;
assign testcases[460] = 64'h8fefbb75110282f0;
assign testcases[461] = 64'h7dcfff9e4b976200;
assign testcases[462] = 64'hdf5eacffdbd79200;
assign testcases[463] = 64'hfdcf9cfefbb66200;
assign testcases[464] = 64'h5c8fffc871c0660d;
assign testcases[465] = 64'hebcf5c96700387fb;
assign testcases[466] = 64'h5f1b06b6f8bb6520;
assign testcases[467] = 64'h0e5fcea780d2f596;
assign testcases[468] = 64'hffef8c3711808506;
assign testcases[469] = 64'hfbcf6edcf8f28000;
assign testcases[470] = 64'h6770d2fadf6e1800;
assign testcases[471] = 64'haf5c383390f38401;
assign testcases[472] = 64'hfd990a4fdffac560;
assign testcases[473] = 64'hfa770a4fdffae460;
assign testcases[474] = 64'h0e5ffdf6a04216f7;
assign testcases[475] = 64'hff9c470250f3d614;
assign testcases[476] = 64'hfc9f3b0460f2f98e;
assign testcases[477] = 64'h7d6fdfa7410081f0;
assign testcases[478] = 64'h4f0a11a0f7cf2d04;
assign testcases[479] = 64'h6b9ffeb8530080f0;
assign testcases[480] = 64'h7effff6d59c59002;
assign testcases[481] = 64'hffbf6b2703409324;
assign testcases[482] = 64'h0f8ffec8a17004f4;
assign testcases[483] = 64'hff8d3823a0f37502;
assign testcases[484] = 64'h1f9af5c0240a0fef;
assign testcases[485] = 64'h4e080280f5fbbf2f;
assign testcases[486] = 64'h3e0a3480e2f8de7f;
assign testcases[487] = 64'h290360d3f9ef8f4a;
assign testcases[488] = 64'hb7ec8f0d18c9f5e0;
assign testcases[489] = 64'h5f5ba780033a7fff;
assign testcases[490] = 64'h7ffffc96401307d5;
assign testcases[491] = 64'hff8c06c6faefd7c0;
assign testcases[492] = 64'h4c5fefabc9f49000;
assign testcases[493] = 64'h0c1f6f49152191f0;
assign testcases[494] = 64'h096daf9a842050f0;
assign testcases[495] = 64'h0a8dfffecab794b0;
assign testcases[496] = 64'h0e18d9d140084fff;
assign testcases[497] = 64'h0c1fbfca851150f0;
assign testcases[498] = 64'h0e7fffec99c59210;
assign testcases[499] = 64'h8d79420056bbffad;
assign testcases[500] = 64'hffbf5f3a8aa35000;
assign testcases[501] = 64'h0288de4f5af6d012;
assign testcases[502] = 64'h0f8ffed7b19075f5;
assign testcases[503] = 64'h7f0b0370e4fbaf2d;
assign testcases[504] = 64'h0e9ffdd6802135c6;
assign testcases[505] = 64'h2e099ac340296fff;
assign testcases[506] = 64'h5f1baab400073fff;
assign testcases[507] = 64'h7bc6900287fbdf4d;
assign testcases[508] = 64'h5c5effed9a672300;
assign testcases[509] = 64'h1f0d59f9ffcca670;
assign testcases[510] = 64'hbf8d280896f8f6e0;
assign testcases[511] = 64'hfb9f0c87f16087fc;
assign testcases[512] = 64'h0e6fffeb973450f0;
assign testcases[513] = 64'hff9f1f0a78c47021;
assign testcases[514] = 64'h0d6fdde6b05477f8;
assign testcases[515] = 64'h5cefffdcd7b30000;
assign testcases[516] = 64'h5f0d08a8fce9d4c0;
assign testcases[517] = 64'h0c6fac85211281f0;
assign testcases[518] = 64'h2f3bd6c00278fd5f;
assign testcases[519] = 64'h199cffefac682400;
assign testcases[520] = 64'h2c7f5c4671f08100;
assign testcases[521] = 64'h4e0ca8c210175dff;
assign testcases[522] = 64'h0a3f4d46112090f1;
assign testcases[523] = 64'h0e8fab85602586f6;
assign testcases[524] = 64'h49deffeae37000f0;
assign testcases[525] = 64'h7f2d0731a0f3fa9b;
assign testcases[526] = 64'h4c9fbb86310182f0;
assign testcases[527] = 64'h6acf2e57b00148fc;
assign testcases[528] = 64'h7d7c8f77600282f2;
assign testcases[529] = 64'h3e08c9a100182fff;
assign testcases[530] = 64'h1ffffca7611004e4;
assign testcases[531] = 64'h1f0d18d9fceae5e0;
assign testcases[532] = 64'h2d199540140a6fff;
assign testcases[533] = 64'hbf4c0710a0f59622;
assign testcases[534] = 64'h4d9fcc97430281f0;
assign testcases[535] = 64'h8fdffdc9d6e28001;
assign testcases[536] = 64'h0f7fffaa550006c6;
assign testcases[537] = 64'hff6f0a646066ecef;
assign testcases[538] = 64'hcb5f2be7f110069c;
assign testcases[539] = 64'h6f0c0540b1f6fc8b;
assign testcases[540] = 64'h1f0c0956b9b7b3f0;
assign testcases[541] = 64'h3e09a9b2202a5fff;
assign testcases[542] = 64'h0c6fdcb6901466f6;
assign testcases[543] = 64'h0f9ffdd7a16074f5;
assign testcases[544] = 64'h9e5f1a0470f38530;
assign testcases[545] = 64'h5f1b0460e3f9be3f;
assign testcases[546] = 64'h3f0d0a16f5d7b3f0;
assign testcases[547] = 64'hde5d0720b3f9ff8d;
assign testcases[548] = 64'h9e4be6d015aaff0f;
assign testcases[549] = 64'h0f2f9ffefab77440;
assign testcases[550] = 64'h0d7ffef8d2a074f4;
assign testcases[551] = 64'h0f3f3b2674e7f5f0;
assign testcases[552] = 64'h098cfffcb78340f1;
assign testcases[553] = 64'h7cbffec9550383f0;
assign testcases[554] = 64'h5d98b250260b8eff;
assign testcases[555] = 64'h0fdffdfaf8d59290;
assign testcases[556] = 64'h0f8fcc98540080f1;
assign testcases[557] = 64'h1a3f9f78130180f0;
assign testcases[558] = 64'hd8ffafcaf9d17001;
assign testcases[559] = 64'haf3e0897fada6510;
assign testcases[560] = 64'hcf0f3a9480157aff;
assign testcases[561] = 64'h3c7fbd88f7f28001;
assign testcases[562] = 64'h4dacbf0ecdf8a410;
assign testcases[563] = 64'h7caffec8720080f0;
assign testcases[564] = 64'h2f3bb5c00378fc6f;
assign testcases[565] = 64'h6e2951c0f6ee7f0d;
assign testcases[566] = 64'h7d9fffebb7e37100;
assign testcases[567] = 64'h2e8fdc88e6f28000;
assign testcases[568] = 64'hffae5a2602609424;
assign testcases[569] = 64'h8e8f0b47f8fca660;
assign testcases[570] = 64'h7f4c0845d7f8c490;
assign testcases[571] = 64'hff6f0903b2f64530;
assign testcases[572] = 64'h0d6ad5a075dbff4e;
assign testcases[573] = 64'hffad592470d36401;
assign testcases[574] = 64'h3f9f9b560230a0f0;
assign testcases[575] = 64'h9b8f1b86a00248fc;
assign testcases[576] = 64'h7f2ba77000287fff;
assign testcases[577] = 64'h5a6f9b750354b0f4;
assign testcases[578] = 64'h1d6fab650234a2f0;
assign testcases[579] = 64'h7f1ad7a100274eff;
assign testcases[580] = 64'hff8f3a0460f2b614;
assign testcases[581] = 64'h5edfdc68f6f17003;
assign testcases[582] = 64'h36b57044b9ff8f0c;
assign testcases[583] = 64'h6cc9f36066dbef0d;
assign testcases[584] = 64'hcf0ebaf45015aaff;
assign testcases[585] = 64'haf3f9dbff9f28003;
assign testcases[586] = 64'h4c4f8b750281f0f5;
assign testcases[587] = 64'h6e4670e2f9df6f0c;
assign testcases[588] = 64'hee4f08714048fdcf;
assign testcases[589] = 64'haccffd99f8f39000;
assign testcases[590] = 64'hffaf3c8ceea86300;
assign testcases[591] = 64'hac4f0bb6e0449aff;
assign testcases[592] = 64'h4f5f0a47f7fab580;
assign testcases[593] = 64'h3d6ad5d064095eff;
assign testcases[594] = 64'h097cefffecc8c4d0;
assign testcases[595] = 64'h6d1e0640c1f8ef7f;
assign testcases[596] = 64'h3f6f0c08a9f8c4b0;
assign testcases[597] = 64'h8c3b0180f6ff8f0b;
assign testcases[598] = 64'hfeaf3c47c8e26004;
assign testcases[599] = 64'h3d8fbd88f6f18001;
assign testcases[600] = 64'hbf5c280430c0f474;
assign testcases[601] = 64'hee8c0c5fdfeae5f0;
assign testcases[602] = 64'hcf6c0879fafbd6c0;
assign testcases[603] = 64'h0d3faf9a763290f0;
assign testcases[604] = 64'hff6f6ab550046aaf;
assign testcases[605] = 64'h5e2d0640c0f7de5f;
assign testcases[606] = 64'h2e09a67023295fff;
assign testcases[607] = 64'hff4c09f9fedb6610;
assign testcases[608] = 64'h9f6f2b0641f0f471;
assign testcases[609] = 64'h09dbff1e38b30065;
assign testcases[610] = 64'h0b6ccefffcf8e4e0;
assign testcases[611] = 64'h5f0a66f7edbea780;
assign testcases[612] = 64'h2b7f8c76300080f0;
assign testcases[613] = 64'h0a4baeffecb88470;
assign testcases[614] = 64'h9dfffdd9d4b000c0;
assign testcases[615] = 64'h3d69fe5f8bf9c100;
assign testcases[616] = 64'hdf6cf6f00067fd6f;
assign testcases[617] = 64'h1f19a890330b6fff;
assign testcases[618] = 64'h1e8ffda9f8f38002;
assign testcases[619] = 64'h3c8fab76200281f0;
assign testcases[620] = 64'h0d6fdc69b8f3a022;
assign testcases[621] = 64'h2e8fac58050180f0;
assign testcases[622] = 64'h3fafa982500686f6;
assign testcases[623] = 64'h3c56201498fd9f0e;
assign testcases[624] = 64'h3f0c07a7fafbf5f0;
assign testcases[625] = 64'hffaebaffeac47100;
assign testcases[626] = 64'h96faff8d76900126;
assign testcases[627] = 64'h0b2490f4fc9f1e16;
assign testcases[628] = 64'h3d6fce7ac8f49100;
assign testcases[629] = 64'h6d689220052b8fff;
assign testcases[630] = 64'hca9f0ca6f02279fe;
assign testcases[631] = 64'h0a5ddffeebd7c4d0;
assign testcases[632] = 64'h0f6fcffcf6f0b2c5;
assign testcases[633] = 64'h0720a1f6feaf4a23;
assign testcases[634] = 64'h0b5fcf6aa6f28002;
assign testcases[635] = 64'h2c069770322a6fff;
assign testcases[636] = 64'h2dbfed89c8f4a000;
assign testcases[637] = 64'h0e4fbdc7b19084f4;
assign testcases[638] = 64'h4fff8f0c39e7b200;
assign testcases[639] = 64'hdf6f0b0470f2a420;
assign testcases[640] = 64'hfcdf1e2aecf8b300;
assign testcases[641] = 64'h3e3690f4fc8f0c05;
assign testcases[642] = 64'h9fffaf4b88d58100;
assign testcases[643] = 64'h4fbffd9af6f28002;
assign testcases[644] = 64'hfe8d3f9faab47003;
assign testcases[645] = 64'h9edfdda9f8c46200;
assign testcases[646] = 64'hbfffee8c58956100;
assign testcases[647] = 64'h0faffde8b38055e6;
assign testcases[648] = 64'h9daffeead6c26000;
assign testcases[649] = 64'h6b9ffdd7720072f0;
assign testcases[650] = 64'h1fcf6a0fbff7b011;
assign testcases[651] = 64'h075abdfffdd8b4a0;
assign testcases[652] = 64'h9f7f0c8afdca8550;
assign testcases[653] = 64'hffad693511808302;
assign testcases[654] = 64'h0d6fbfa79063a5f5;
assign testcases[655] = 64'h08197deffec99580;
assign testcases[656] = 64'h9fdfdc79f7f28000;
assign testcases[657] = 64'h3c0fcffcc6c0f546;
assign testcases[658] = 64'h8f1e29f8fdb96400;
assign testcases[659] = 64'hffaf5b1611909302;
assign testcases[660] = 64'hff8d290440e1a403;
assign testcases[661] = 64'h6f0c09eafc8d4710;
assign testcases[662] = 64'hff9c4722a0f38503;
assign testcases[663] = 64'h0f5fad792642a1f0;
assign testcases[664] = 64'h6aaffde6720073f0;
assign testcases[665] = 64'h0d2f9fffecb88460;
assign testcases[666] = 64'hfd4f0e0b283543a0;
assign testcases[667] = 64'h6fef5f29a8f48003;
assign testcases[668] = 64'h8fcfecbaf6d27001;
assign testcases[669] = 64'h4e9feeebf7e48100;
assign testcases[670] = 64'haf3c0630c0f59816;
assign testcases[671] = 64'h0b6cffffcca894d0;
assign testcases[672] = 64'hffffdcaa87652200;
assign testcases[673] = 64'haf59fbcf9af9b001;
assign testcases[674] = 64'h785fdfe8830070f0;
assign testcases[675] = 64'hacefcda8720081f1;
assign testcases[676] = 64'h3d0650d1f8ce4f0a;
assign testcases[677] = 64'h8f1f7daef9f39001;
assign testcases[678] = 64'h1730b0f6dc6f1a04;
assign testcases[679] = 64'hdf2d86f05089bf0b;
assign testcases[680] = 64'hef8c371290f28402;
assign testcases[681] = 64'heb8f0c76c03399fe;
assign testcases[682] = 64'h0c6fdfebb7f3a043;
assign testcases[683] = 64'h2e5f8c570333a3f0;
assign testcases[684] = 64'h0f28c880220b6fff;
assign testcases[685] = 64'h299dffdca7820030;
assign testcases[686] = 64'h4eafb963002593f3;
assign testcases[687] = 64'h6ccfcda5600181f1;
assign testcases[688] = 64'hfc9f0d38dbebd5d0;
assign testcases[689] = 64'h4f6bfe4f0dcac550;
assign testcases[690] = 64'h0b0560e1f7cd5f1b;
assign testcases[691] = 64'hbffffbb8f4c06001;
assign testcases[692] = 64'h7c4bf6c074faff0d;
assign testcases[693] = 64'h0072d5faef6f4cba;
assign testcases[694] = 64'h6fffff6f8bf6a100;
assign testcases[695] = 64'h0d1f9fffecc8b490;
assign testcases[696] = 64'hbf4b061090f4faef;
assign testcases[697] = 64'h4ebfdca8540080f0;
assign testcases[698] = 64'h086abdfffce8d4f0;
assign testcases[699] = 64'hff9e3a0450d2a614;
assign testcases[700] = 64'h9aaffdd680e39809;
assign testcases[701] = 64'h4d6fcc88b8f39002;
assign testcases[702] = 64'haf0f4a74000599fe;
assign testcases[703] = 64'h0d5fce6b88f6b230;
assign testcases[704] = 64'h4831a0f5fd9f1d06;
assign testcases[705] = 64'hfe8f5a9410058aff;
assign testcases[706] = 64'h3daffda9c7f49100;
assign testcases[707] = 64'h3b0450c2f8ce5f0c;
assign testcases[708] = 64'h0fbffcc8836004b5;
assign testcases[709] = 64'h5fef7f1b9af6a200;
assign testcases[710] = 64'h3f498440160c7fff;
assign testcases[711] = 64'h5d8ffed8640493f0;
assign testcases[712] = 64'h1b4fcfaa560170f1;
assign testcases[713] = 64'h7fffda85200548f8;
assign testcases[714] = 64'h8b0b85e04289ff7e;
assign testcases[715] = 64'hccdf1f09b9fbc590;
assign testcases[716] = 64'haeeffde9e4a15002;
assign testcases[717] = 64'h88290081e8ff8d17;
assign testcases[718] = 64'h1e8fff9bc8f58200;
assign testcases[719] = 64'h072abdffcca88460;
assign testcases[720] = 64'hbf7cb570041b7fff;
assign testcases[721] = 64'h5dafecb7630081f2;
assign testcases[722] = 64'h8f1bfabf4900e127;
assign testcases[723] = 64'hff8c380440f1c405;
assign testcases[724] = 64'hff9e3a0430b2a737;
assign testcases[725] = 64'h1f2f0a0594e7e5f0;
assign testcases[726] = 64'hff9e5a2540e1b507;
assign testcases[727] = 64'h5c8fdcb6520080f0;
assign testcases[728] = 64'h5f191390f4faaf0f;
assign testcases[729] = 64'h3b9fffcb97f49001;
assign testcases[730] = 64'hff0cf9dfa701f088;
assign testcases[731] = 64'h078cffdcb7a10050;
assign testcases[732] = 64'h0e7ffcd6908116d6;
assign testcases[733] = 64'hbf4d180440f0f471;
assign testcases[734] = 64'h3eafbb660220a0f0;
assign testcases[735] = 64'h0d2f3c3844b3e4f0;
assign testcases[736] = 64'h2f196310081f8fff;
assign testcases[737] = 64'h0d5fbf99451180f0;
assign testcases[738] = 64'haf0dabf580156b7f;
assign testcases[739] = 64'h0548acffdd986440;
assign testcases[740] = 64'h4f6cb670250c5fff;
assign testcases[741] = 64'h5fefdf5c89f59003;
assign testcases[742] = 64'h3f3ba650030c7fff;
assign testcases[743] = 64'h0f8ffed9a4703597;
assign testcases[744] = 64'h5cbfcf9a843000f0;
assign testcases[745] = 64'h9bcfab84500080f1;
assign testcases[746] = 64'h5ebfffdbb8b46100;
assign testcases[747] = 64'h5f0c9d7cc8f4c021;
assign testcases[748] = 64'h0e5f7c470351a0f0;
assign testcases[749] = 64'h4fafcc79f7f38001;
assign testcases[750] = 64'h5effffaa550015b6;
assign testcases[751] = 64'h8b7f1c96800379fe;
assign testcases[752] = 64'h3e090360d4f9df6f;
assign testcases[753] = 64'hcf8b640057bcff7c;
assign testcases[754] = 64'h0c8effcdaa764310;
assign testcases[755] = 64'h4fffdf4c8af7b100;
assign testcases[756] = 64'h2f2ac7a001095fff;
assign testcases[757] = 64'haccffcc7820080f1;
assign testcases[758] = 64'hff8f1c0742e0f464;
assign testcases[759] = 64'h5b9fecb6420282f0;
assign testcases[760] = 64'hff3d76a00279cf0c;
assign testcases[761] = 64'h7fefcc98f5e07003;
assign testcases[762] = 64'hff9d593460d08301;
assign testcases[763] = 64'h0c5fbe98440081f0;
assign testcases[764] = 64'h8f1db7f013c9ff0e;
assign testcases[765] = 64'hee5a0e9febf5f031;
assign testcases[766] = 64'h1f3c0676f5cbc4d0;
assign testcases[767] = 64'h0a7cdffffce7c3e0;
assign testcases[768] = 64'h0fbfedc6a06237f8;
assign testcases[769] = 64'h0e5fbd88343090f0;
assign testcases[770] = 64'h5c0710a2f8fe7f1b;
assign testcases[771] = 64'h7f2b0450c1f7ed7f;
assign testcases[772] = 64'hff9e49051091a514;
assign testcases[773] = 64'hfc8f0d87b0044bff;
assign testcases[774] = 64'hfd8f0e3acbf8c240;
assign testcases[775] = 64'h0668ccffdda97440;
assign testcases[776] = 64'hff9f5d99e5d16000;
assign testcases[777] = 64'h0f498410161d7fff;
assign testcases[778] = 64'hcc8f0ca7f04057fc;
assign testcases[779] = 64'h4c7fab750262d0f5;
assign testcases[780] = 64'h6cd7f081c8fe9f0c;
assign testcases[781] = 64'h089cfffee8e370f1;
assign testcases[782] = 64'h04a7fe8f59e49014;
assign testcases[783] = 64'hde9cadafc9e200f0;
assign testcases[784] = 64'h6f4f0740d2f9af3c;
assign testcases[785] = 64'hff9d5843a0f48603;
assign testcases[786] = 64'h8fae4a0695f9d4c0;
assign testcases[787] = 64'h2e9fbc89f7f28002;
assign testcases[788] = 64'hffaf3e1878c58100;
assign testcases[789] = 64'h0f7fbca6804596f6;
assign testcases[790] = 64'hcf7c280390f48714;
assign testcases[791] = 64'h0eafecb6704065f6;
assign testcases[792] = 64'h0b7dfffedaa76340;
assign testcases[793] = 64'h0a6dcfffcb884440;
assign testcases[794] = 64'hcefffca9e6d27000;
assign testcases[795] = 64'h0f5ffdd790f1d617;
assign testcases[796] = 64'h9deffc89f6f28002;
assign testcases[797] = 64'h1c6fee89d8f39002;
assign testcases[798] = 64'h3fbffd890623c2f0;
assign testcases[799] = 64'haf6f5c9ed8f3a001;
assign testcases[800] = 64'hff8f2a0290f46611;
assign testcases[801] = 64'h0d69e6b022094eff;
assign testcases[802] = 64'h41a8ff8f49d5b000;
assign testcases[803] = 64'h4ea9f330059aff4f;
assign testcases[804] = 64'h6f1a0380f4fabf3e;
assign testcases[805] = 64'hff8f2d1788d48001;
assign testcases[806] = 64'h0558acfffde9c4b0;
assign testcases[807] = 64'h9f1b888000277eff;
assign testcases[808] = 64'h7de7f03005aaef1f;
assign testcases[809] = 64'h8a8fffe8820081f0;
assign testcases[810] = 64'hbf7f291380f38502;
assign testcases[811] = 64'h6b8f6c66410081f2;
assign testcases[812] = 64'h7faf9a550251a0f0;
assign testcases[813] = 64'hde7f1b0540c2f7ee;
assign testcases[814] = 64'h2c6fac87420080f0;
assign testcases[815] = 64'h8d8fffcbc8f37001;
assign testcases[816] = 64'h7e7fef9ab9f4a000;
assign testcases[817] = 64'h2f1b2b0d350031f2;
assign testcases[818] = 64'h098cffefebe8e4d0;
assign testcases[819] = 64'h9cbffcc8640060f0;
assign testcases[820] = 64'h7f1c0796f7cc9660;
assign testcases[821] = 64'h1f3f09a6f9de8750;
assign testcases[822] = 64'h4f0b0370e3facf5f;
assign testcases[823] = 64'h0a4f9c85302294f2;
assign testcases[824] = 64'h0a5bbefffcd8b4a0;
assign testcases[825] = 64'h8bc6f08177ccaf0d;
assign testcases[826] = 64'hffae592380f46401;
assign testcases[827] = 64'h3f18a870030d7fff;
assign testcases[828] = 64'h6bdb8f0746b0f824;
assign testcases[829] = 64'h2c6fee9af7f27001;
assign testcases[830] = 64'h5f3c0814c6e8e4f0;
assign testcases[831] = 64'h8fffef4e9af5a000;
assign testcases[832] = 64'h097dcfbaa55051f1;
assign testcases[833] = 64'h5f4ba550043b7fff;
assign testcases[834] = 64'h0f8efca6402265f6;
assign testcases[835] = 64'hde6f4acdfdf79100;
assign testcases[836] = 64'h0e8fffccc8e58200;
assign testcases[837] = 64'hdf8d4834b2f57300;
assign testcases[838] = 64'h2c8fbf89620180f0;
assign testcases[839] = 64'h1f38f8b010093fff;
assign testcases[840] = 64'hff9f3b0530b09422;
assign testcases[841] = 64'hff8d390520b0a321;
assign testcases[842] = 64'h290731b0f5fcaf3f;
assign testcases[843] = 64'h5f099890312a7fff;
assign testcases[844] = 64'hcf6d282390f3a708;
assign testcases[845] = 64'h0c6fdeb7612093f0;
assign testcases[846] = 64'haf6d290494f7b490;
assign testcases[847] = 64'h5f2c0886f9f9d4a0;
assign testcases[848] = 64'h6f2c0766f6f8e4b0;
assign testcases[849] = 64'h0c7f8f7872f1b050;
assign testcases[850] = 64'hff0f49e28046fc6f;
assign testcases[851] = 64'h0f8fffc9a27084f3;
assign testcases[852] = 64'h0f8fddb7905477f8;
assign testcases[853] = 64'h6f8b07a6f6ead5c0;
assign testcases[854] = 64'h5e0a0380f4fbbf4c;
assign testcases[855] = 64'h8f397c8d740060f0;
assign testcases[856] = 64'h0b9dcffefaf7d3e0;
assign testcases[857] = 64'h3f0a0460e3f9cf5d;
assign testcases[858] = 64'h0f7feffdba967320;
assign testcases[859] = 64'h0b3f9f89540090f1;
assign testcases[860] = 64'h5e9f9a560241a1f0;
assign testcases[861] = 64'hdd9f3daaf8f38000;
assign testcases[862] = 64'h8deffbd6810080f0;
assign testcases[863] = 64'h4b8fcc86120281f0;
assign testcases[864] = 64'had280092f8ff7f09;
assign testcases[865] = 64'h0f6fad9ab6f4c160;
assign testcases[866] = 64'h0faffde8d3b064f6;
assign testcases[867] = 64'h7d4fac66020080f0;
assign testcases[868] = 64'hfe8f4b75600358cb;
assign testcases[869] = 64'hbf8afd9fece89001;
assign testcases[870] = 64'h5f2c0796f7cb9670;
assign testcases[871] = 64'haf4d080380f3a634;
assign testcases[872] = 64'haffcffacfdf5b001;
assign testcases[873] = 64'h5bafaf9a740030f0;
assign testcases[874] = 64'h0779ccffdca87460;
assign testcases[875] = 64'h0f4afd6f99f7c024;
assign testcases[876] = 64'hef2f49f480047aff;
assign testcases[877] = 64'h0e097540140b7fff;
assign testcases[878] = 64'h082a9dfffcc89450;
assign testcases[879] = 64'h4f2c06a5fafbe6c0;
assign testcases[880] = 64'h8f2d0630a0f4faac;
assign testcases[881] = 64'h7b9ffdc8630081f0;
assign testcases[882] = 64'h0a6defffecc8b4b0;
assign testcases[883] = 64'hff9f6cfdecb87300;
assign testcases[884] = 64'h0d4fdfdcd8f49200;
assign testcases[885] = 64'h4ebffdcad6f28000;
assign testcases[886] = 64'h0c5f9b76211393f0;
assign testcases[887] = 64'hcdfffdd9b6b15001;
assign testcases[888] = 64'h6f3c0896f8d9a470;
assign testcases[889] = 64'h0e7feec7a06377f8;
assign testcases[890] = 64'h4fbfaa65010280f0;
assign testcases[891] = 64'hf8680b4fcfe9c450;
assign testcases[892] = 64'h1d8fffba77e48001;
assign testcases[893] = 64'hef8d07c7fbeec7a0;
assign testcases[894] = 64'h3f1841b0f6ed7f0d;
assign testcases[895] = 64'h4d1650d2f9cf4f08;
assign testcases[896] = 64'h0e6fefb8805386f8;
assign testcases[897] = 64'h5ecfdc78e7f39000;
assign testcases[898] = 64'h0d7fffea972340f0;
assign testcases[899] = 64'h2b4f7c450042a1f0;
assign testcases[900] = 64'hbe19fc7f5700e224;
assign testcases[901] = 64'hafffef8db9d37002;
assign testcases[902] = 64'hfe5f7af46005caff;
assign testcases[903] = 64'h0a7defffdcb89470;
assign testcases[904] = 64'h6f0a33e2f6cea890;
assign testcases[905] = 64'h9e3e0740c2f9df6f;
assign testcases[906] = 64'h3f2b1652e2f47300;
assign testcases[907] = 64'h6f3a04d4f8ceb7b0;
assign testcases[908] = 64'h9ccffbb5420382f0;
assign testcases[909] = 64'h0c2f9faa652090f1;
assign testcases[910] = 64'h0f9fcd97804376f6;
assign testcases[911] = 64'h5f3d0825c6f9e4e0;
assign testcases[912] = 64'h5f6a9330062d9ffd;
assign testcases[913] = 64'h8fffacbaf6d26001;
assign testcases[914] = 64'h0faffcd7927045f6;
assign testcases[915] = 64'h0b4fcfc8928085f6;
assign testcases[916] = 64'h1d7f9b66020181f0;
assign testcases[917] = 64'hcf4f6ab440057aff;
assign testcases[918] = 64'h084abeffcc884420;
assign testcases[919] = 64'h5b9fcc96510180f0;
assign testcases[920] = 64'h6caf9b660544a1f0;
assign testcases[921] = 64'hdf0e0adcffdbb590;
assign testcases[922] = 64'h0e4f9e784350b0f2;
assign testcases[923] = 64'h6f1c0673e5f9b580;
assign testcases[924] = 64'h5eafcb67032190f0;
assign testcases[925] = 64'h0c6fac96604266f7;
assign testcases[926] = 64'h2f0c8950041e7fff;
assign testcases[927] = 64'hfc7c6ffffbd77300;
assign testcases[928] = 64'h7ecfdba8f5c16001;
assign testcases[929] = 64'hfc9f0c88ecf6d010;
assign testcases[930] = 64'h7cafffcb670340d0;
assign testcases[931] = 64'h5c180350d2f6fbdf;
assign testcases[932] = 64'hbf5b0540c3f9ef5f;
assign testcases[933] = 64'h7d3a8420042b7fff;
assign testcases[934] = 64'h5840f0ca662fbf0c;
assign testcases[935] = 64'h4f2c0785f6dab5b0;
assign testcases[936] = 64'h0c4f8e692442a1f0;
assign testcases[937] = 64'h5f7ae6a002294fff;
assign testcases[938] = 64'h5f3c07b5faeb9540;
assign testcases[939] = 64'h0f8ffeea87f4b130;
assign testcases[940] = 64'h1d0640c2f8df6f1a;
assign testcases[941] = 64'h5e69af0a4760f748;
assign testcases[942] = 64'hbf0e47d00077fe3f;
assign testcases[943] = 64'h08299dfffcb88450;
assign testcases[944] = 64'h4d9fcb95320181f0;
assign testcases[945] = 64'h0a2a8deffde8c490;
assign testcases[946] = 64'h2f9f9c58050281f0;
assign testcases[947] = 64'h6e598320069bff3f;
assign testcases[948] = 64'h9fabe580240c6fff;
assign testcases[949] = 64'h4c5fac66011080f1;
assign testcases[950] = 64'h4e1a9740130b6fff;
assign testcases[951] = 64'h0f8fffd9b29075f7;
assign testcases[952] = 64'h0f4fbfb8a07185f3;
assign testcases[953] = 64'hae3a0450c4facf4f;
assign testcases[954] = 64'h2e5fffca76f3a001;
assign testcases[955] = 64'hbbff6f0c8cc98430;
assign testcases[956] = 64'h1c5fdfbbf7f28001;
assign testcases[957] = 64'h5f2e0a89fca96430;
assign testcases[958] = 64'hfe4f0bbbffebc5b0;
assign testcases[959] = 64'h2b9ffca6500255f5;
assign testcases[960] = 64'h1f3d0824b4f8f5e0;
assign testcases[961] = 64'h0b0a48a420285fff;
assign testcases[962] = 64'hff9e3a0501809403;
assign testcases[963] = 64'h0d7ddffffce8c4c0;
assign testcases[964] = 64'h0f5fcf98403176f8;
assign testcases[965] = 64'h3f1d08a7fbe9b580;
assign testcases[966] = 64'h2d0560d3fbaf3b24;
assign testcases[967] = 64'h9f0f4caeebf5a000;
assign testcases[968] = 64'hbe0f38d22076fc8f;
assign testcases[969] = 64'h4c6ffffcb8f48100;
assign testcases[970] = 64'hcbaf0c96d00268fe;
assign testcases[971] = 64'h4f096980303b7fff;
assign testcases[972] = 64'hef6d07b6f9ceb7b0;
assign testcases[973] = 64'h0fffdba6803014f6;
assign testcases[974] = 64'h9dffef6c47b58100;
assign testcases[975] = 64'h5f0e17e7fdbfb8c0;
assign testcases[976] = 64'h5d080190f5fc8f1c;
assign testcases[977] = 64'h1e7f9b56022190f0;
assign testcases[978] = 64'h0f1cb6f07188de4f;
assign testcases[979] = 64'hffbf6b2702608406;
assign testcases[980] = 64'h06488acdffdcb6a0;
assign testcases[981] = 64'h7dafdc88f7f37001;
assign testcases[982] = 64'hff8f2a0450e2c718;
assign testcases[983] = 64'h4e69fc4f7df8d200;
assign testcases[984] = 64'h7f3d0835a5f6e4d0;
assign testcases[985] = 64'heeffaf9bd6c16000;
assign testcases[986] = 64'h4a945003a7fd8f0c;
assign testcases[987] = 64'hff9f4b0530b3f8ee;
assign testcases[988] = 64'h4e0aa79000185fff;
assign testcases[989] = 64'hff9f2c0722a0c447;
assign testcases[990] = 64'h5b3a3400077cff7f;
assign testcases[991] = 64'h55086cfffdd8c4c0;
assign testcases[992] = 64'h6d9fecb7530493f0;
assign testcases[993] = 64'hffae4a0601708425;
assign testcases[994] = 64'hcf7b4620b0f47502;
assign testcases[995] = 64'h3f3b5f78a10051f2;
assign testcases[996] = 64'h4eafacb8f5d17000;
assign testcases[997] = 64'h1f2ba650041c5fff;
assign testcases[998] = 64'h9d1f2ae5b00499ff;
assign testcases[999] = 64'h8d9fffd8730072f0;


  
  localparam SUM_BITS = $clog2(HIDDEN_CNT+1);
  wire [$clog2(CLASS_CNT)-1:0] prediction;

  // Instantiate module under test
 pendigits_ts #(
 ) dut (
    .data(data),
    .clk(clk),
    .rst(rst),
    .prediction(prediction)
  );
  
  always #halfT clk <= ~clk;

  integer i;
  initial begin
    $write("["); //" 
    for(i=0;i<TEST_CNT;i=i+1)
        runtestcase(i);
    $display("]");
    $finish;
  end

  task runtestcase(input integer i); begin
    data <= testcases[i];
    rst <= 1;
    clk <= 0;
    #period
    rst <= 0;
    #period
    #((FEAT_CNT+HIDDEN_CNT-1)*period)
    $write("%d, ",prediction);
  end
  endtask

endmodule
