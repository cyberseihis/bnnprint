












module gasId_bnn1_bnnseq #(

parameter FEAT_CNT = 128,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 6,
parameter TEST_CNT = 1000


  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] features,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  localparam Weights0 = 5120'b10101110011001110100010101110101000111001100101001000001000110101111111111000010010010110011001110100001111101011101010110001011000001110010000111110101010001001000100101000001101010101111110101001101110011000000111010011000110000101111000000100110100100011010010000110111011000100011000110010011001011110011110011010100101111110110001100010011010111011101110010111111010000011000000101011001110101011010110100101111000000000111010111010100100010010010111111100110011111011101010010101101111000111001001100011111110111000001001001110110101110111101000000001101101111010011101111000011000110000111101100001010100101101001000011111111001000110111010111000010110110111000111110010010011101111111100010111100100100100101000101111101111110001111111010101010101000110111000011100000100010001001001111000101011011001100010000100010111011010010011011011110000010110001011010100111010010101100110010000010111001100101000011010100110110111010101010111011101111111111111111110101010110100101010000011110110000100111001011111000101111101001101000111111011101011111000011111100000010101001000101110001111110001011110011110010001011011101111000000111010110010011010100111010010111000000110111110000110101110100011011000101111000010001001001010011100010000000000100010110100010010001101101111100000111010101011101001101100010101001000010000101111101010000011111111001110111011001110001011111111001110110011000100010110110100100001000011011101101010010011110010101111101111111011001000001110110010110011110110001010101000011101011110011001011011000111011111011101011011011100111110010101100001110011110011011100110101001010000001000011111010000111010101010111100110000100111110110010111010010111110001001000101101110010101100110001000101101101001000010000110111010010100100011010111011011100000110100010010100111110100101101011010000011011010110100010101000011101010111100101011111110010001010110011110001101100111101101001001000111010011110011101100110111010100000101100101011111100100000111101011101111011110111100001001110101101100001000000100100010001111110010110010000011111010110001001000110101101000000010000010111001010100100111110010000110010111011010000101010000101111000111100110101011101101100001001111000001000011011101001011010010100101011010011001011110101011100111000111011000000010011111000111100111100101010111011010001110100011000001010110010111010001100110010010001101100000011101110101000010011100011010110110010110100111110101001001100001010011001110100011001001101111000001011001011110101000000001111110100000101100110111001111110000011101100000111000001010101000100011000000111111010111010100100010000011111101100110011101000110110010101110001001110000000101111101000101101000101000100111000000110111010101011100100111100110001100000011001111011101010000011111111110010110011000111011100101110101101000000111111100010110110110110110001110110000011001100011111110010111111010111010011001110000000110110101000111101000101001001111010011111111010100101110100010100101001100010011011101010001111010001010000001100100001111110101001111101000111001000010000000111001010110010110001110110010101111011011111001111011110010000010001011000011110010001011111100011001100101011111011110111100110110010101111101111111100100010001000111001100110101110101101010000011101010010000010111010011011111101001101001101001001100011101011100101100100000011001100100000010011101010001011000001001000010000000001101011100110100001111001110010010110001101101110110001110010011111001100001110110011100001000101101001010110010000001101011111001010111111011100100110101000111001000011101101111000000111110000110110100010101110101111110111010111000000001001101010100110111010000101110111011000100001111000010000011100011101110111100000110001110110000100001010000101101000101011011111001011001100101010110001110101010100101101000111001001111010010101110001010101011011101110001101100010000000111110110111101000011011100110011100100101001101011010110100100011001111100001001110000001011001010010001100111111111110101001010101101101001000000000110011011010100101111001001000011000011001110010010000000010100100011011101010110010000011101110100111110001111110100011000110010000100111100110111011101001101000001000011101110101011000100100100001110111011000110001010001101110001000111010011010010011010101010110110100100011001001011011101010010011011011010010000000001101110100101001011111011100100100100011101001110000011000100110110001001101101111000110000111010101110111100001011010000000111000011010010110011111011111000100100111001101110011101000110011010100000111101100100000000111100110111011011100011011110110001101001010111101011000000000110011011000100100111010110000101100000011000101100000010111011110111111100110000010101101111000110100110101101101001100110000111010110000101110001010000000110010011000101100010010110101101011110010110000101011000100001110011000101101000001110001001000101010101100100100110101001000011101100000001010101101010010000000001100110110001001011111100101011100010000010111011000101101111010001100001110000001110110011101001100110100110110000101101000001001101000100111111001110011010110100100011001101100000 ;
  localparam Weights1 = 240'b110110100101001100011011001101010010111001110001111110101011111000010000011011011101010111010010111111100000011011101011101110110001111101110111000101000010110010011111011010110001001100011101110111001001101000011111111101110011010001101100 ;

  seq_bnn #(.FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),.Weights0(Weights0),.Weights1(Weights1)) bnn (
    .clk(clk),
    .rst(rst),
    .features(features),
    .prediction(prediction)
  );

endmodule
