











module winewhite_tnn1_tnnzeq #(

parameter FEAT_CNT = 11,
parameter HIDDEN_CNT = 40,
parameter FEAT_BITS = 4,
parameter CLASS_CNT = 7,
parameter TEST_CNT = 1000




  ) (
  input clk,
  input rst,
  input [FEAT_CNT*FEAT_BITS-1:0] data,
  output [$clog2(CLASS_CNT)-1:0] prediction
  );

  seq_tnnzeq #(
      .FEAT_CNT(FEAT_CNT),.FEAT_BITS(FEAT_BITS),.HIDDEN_CNT(HIDDEN_CNT),.CLASS_CNT(CLASS_CNT),
  .SPARSE_VALS(440'b10001100000000000001100000100001001000000010011010001110000011100000010100010000100111101001010000001010111000100001000010000000000001001011000000000000001000000100000001000111101111101101010000011100110000011100001000110000100001000011001110000001000011101111111000001000000010000011100010001010000010100110001010101100000110100010011010000000010001100000000001100011011110000010000001100010100000000100001111000001001101101110000010010000),
  .MASK(440'b10111110001100000001100100111101001011100110011110111110000111111000010100010000100111101001010001101010111010111101011111000000000001001011100100000011001001001101010011101111101111101101010110111111110001011100111100110100111111010111001110001101100111101111111000111001000110110111101010011010011010100110111011101100001110100010111011001011011001111001111001101011011110000110011001100011101100011110011111111101001101101110001110010011),
  .NONZERO_CNT(640'h07030606090603050506090105030508080807070707060904080506080407070707040706080706),
  .SPARSE_VALS2(79'b0100000010110010011000100000110000101111111100111011000110111010101011011001010),  // Bits of not-zeroes
  .COL_INDICES(632'h2625232221201e1b1817141211100d0c0605040201211f17100d0b211c1615100c0825211f1817100f0125242119181412092625221f1e1c1817161413100b0a07261c171412100f0b0a0907060401), // Column of non-zeros
  .ROW_PTRS(64'h4f3a342d251d0e00) // Column of non-zeros // Start indices per row
      ) tnn (
    .clk(clk),
    .rst(rst),
    .features(data),
    .prediction(prediction)
  );

endmodule
